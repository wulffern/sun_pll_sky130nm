magic
tech sky130B
magscale 1 1
timestamp 1720908000
<< checkpaint >>
rect 0 0 3288 2704
<< locali >>
rect 2976 192 3096 2512
rect 192 192 3096 312
rect 192 2392 3096 2512
rect 192 192 312 2512
rect 2976 192 3096 2512
rect 3168 0 3288 2704
rect 0 0 3288 120
rect 0 2584 3288 2704
rect 0 0 120 2704
rect 3168 0 3288 2704
rect 2496 1763 2556 1793
rect 2556 1865 2688 1895
rect 2556 1763 2586 1895
rect 2472 1733 2526 1763
rect 2496 1939 2556 1969
rect 2556 2041 2688 2071
rect 2556 1939 2586 2071
rect 2472 1909 2526 1939
rect 2496 883 2556 913
rect 2556 985 2688 1015
rect 2556 883 2586 1015
rect 2472 853 2526 883
rect 2496 1059 2556 1089
rect 2556 1161 2688 1191
rect 2556 1059 2586 1191
rect 2472 1029 2526 1059
rect 2496 1235 2556 1265
rect 2556 1337 2688 1367
rect 2556 1235 2586 1367
rect 2472 1205 2526 1235
rect 2496 1411 2556 1441
rect 2556 1513 2688 1543
rect 2556 1411 2586 1543
rect 2472 1381 2526 1411
rect 2496 1587 2556 1617
rect 2556 1689 2688 1719
rect 2556 1587 2586 1719
rect 2472 1557 2526 1587
rect 2496 707 2556 737
rect 2556 809 2688 839
rect 2556 707 2586 839
rect 2472 677 2526 707
rect 702 1059 792 1089
rect 600 1337 702 1367
rect 702 1059 732 1367
rect 762 1029 816 1059
<< m3 >>
rect 758 192 866 1088
rect 2850 192 2958 494
rect 2422 192 2530 736
rect 1154 0 1262 1088
rect 2030 2352 2130 2704
rect 2030 2352 2130 2704
rect 2026 384 2134 2704
<< m1 >>
rect 702 531 792 561
rect 600 1161 702 1191
rect 702 531 732 1191
rect 762 501 816 531
rect 762 2674 870 2704
rect 2634 0 2742 30
rect 2634 0 2742 30
rect 2688 457 2772 487
rect 2688 0 2772 30
rect 2772 0 2802 487
rect 762 2674 870 2704
rect 816 1381 900 1411
rect 816 2674 900 2704
rect 900 1381 930 2704
<< m2 >>
rect 600 809 686 847
rect 686 1733 2472 1771
rect 686 809 724 1771
rect 476 457 600 495
rect 476 1909 2472 1947
rect 476 457 514 1947
rect 2472 2085 2558 2123
rect 2558 633 2688 671
rect 2558 633 2596 2123
use SUN_PLL_LSCORE xa3 
transform 1 0 384 0 1 384
box 384 384 1644 1088
use SUNTR_IVX1_CV xa4 ../SUN_TR_SKY130NM
transform 1 0 384 0 1 1088
box 384 1088 1644 1264
use SUNTR_IVX1_CV xa5 ../SUN_TR_SKY130NM
transform 1 0 384 0 1 1264
box 384 1264 1644 1440
use SUNTR_TAPCELLB_CV xa6 ../SUN_TR_SKY130NM
transform 1 0 384 0 1 1440
box 384 1440 1644 1616
use SUNTRB_NDX1_CV xb1 ../SUN_TRB_SKY130NM
transform -1 0 2904 0 1 384
box 2904 384 4164 736
use SUNTRB_IVX1_CV xb2_0 ../SUN_TRB_SKY130NM
transform -1 0 2904 0 1 736
box 2904 736 4164 912
use SUNTRB_IVX1_CV xb2_1 ../SUN_TRB_SKY130NM
transform -1 0 2904 0 1 912
box 2904 912 4164 1088
use SUNTRB_IVX1_CV xb2_2 ../SUN_TRB_SKY130NM
transform -1 0 2904 0 1 1088
box 2904 1088 4164 1264
use SUNTRB_IVX1_CV xb2_3 ../SUN_TRB_SKY130NM
transform -1 0 2904 0 1 1264
box 2904 1264 4164 1440
use SUNTRB_IVX1_CV xb2_4 ../SUN_TRB_SKY130NM
transform -1 0 2904 0 1 1440
box 2904 1440 4164 1616
use SUNTRB_IVX1_CV xb2_5 ../SUN_TRB_SKY130NM
transform -1 0 2904 0 1 1616
box 2904 1616 4164 1792
use SUNTRB_IVX1_CV xb2_6 ../SUN_TRB_SKY130NM
transform -1 0 2904 0 1 1792
box 2904 1792 4164 1968
use SUNTRB_IVX1_CV xb2_7 ../SUN_TRB_SKY130NM
transform -1 0 2904 0 1 1968
box 2904 1968 4164 2144
use SUNTRB_TAPCELLBAVSS_CV xb3 ../SUN_TRB_SKY130NM
transform -1 0 2904 0 1 2144
box 2904 2144 4164 2320
use cut_M1M4_2x1 xcut0 
transform 1 0 762 0 1 192
box 762 192 862 230
use cut_M1M4_2x1 xcut1 
transform 1 0 2854 0 1 192
box 2854 192 2954 230
use cut_M1M4_2x1 xcut2 
transform 1 0 2426 0 1 192
box 2426 192 2526 230
use cut_M1M4_2x1 xcut3 
transform 1 0 1158 0 1 0
box 1158 0 1258 38
use cut_M1M2_2x1 xcut4 
transform 1 0 778 0 1 501
box 778 501 870 535
use cut_M1M2_2x1 xcut5 
transform 1 0 562 0 1 1161
box 562 1161 654 1195
use cut_M1M3_2x1 xcut6 
transform 1 0 546 0 1 809
box 546 809 646 847
use cut_M1M3_2x1 xcut7 
transform 1 0 2418 0 1 1733
box 2418 1733 2518 1771
use cut_M1M3_2x1 xcut8 
transform 1 0 554 0 1 457
box 554 457 654 495
use cut_M1M3_2x1 xcut9 
transform 1 0 2426 0 1 1909
box 2426 1909 2526 1947
use cut_M1M3_2x1 xcut10 
transform 1 0 2418 0 1 2085
box 2418 2085 2518 2123
use cut_M1M3_2x1 xcut11 
transform 1 0 2634 0 1 633
box 2634 633 2734 671
use cut_M1M2_2x1 xcut12 
transform 1 0 2634 0 1 457
box 2634 457 2726 491
use cut_M1M2_2x1 xcut13 
transform 1 0 762 0 1 1381
box 762 1381 854 1415
<< labels >>
flabel locali s 2976 192 3096 2512 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
flabel locali s 3168 0 3288 2704 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel m1 s 762 2674 870 2704 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel m3 s 2030 2352 2130 2704 0 FreeSans 400 0 0 0 VDD_ROSC
port 3 nsew signal bidirectional
flabel m1 s 2634 0 2742 30 0 FreeSans 400 0 0 0 PWRUP_1V8
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 3288 2704
<< end >>
