magic
tech sky130B
magscale 1 2
timestamp 1707433200
<< checkpaint >>
rect 0 0 40552 24888
<< locali >>
rect 40252 0 40552 24888
rect 0 0 40552 300
rect 0 24588 40552 24888
rect 0 0 300 24888
rect 40252 0 40552 24888
rect 300 460 460 572
rect 300 5136 460 5248
rect 4516 8558 5092 8778
rect 4516 3882 5092 4102
<< m3 >>
rect 23120 0 23336 484
rect 39988 404 40328 480
rect 39988 1364 40328 1440
rect 39988 2324 40328 2400
rect 39988 3284 40328 3360
rect 39988 4244 40328 4320
rect 39988 5204 40328 5280
rect 39988 6164 40328 6240
rect 39988 7124 40328 7200
rect 39988 8084 40328 8160
rect 39988 9044 40328 9120
rect 39988 10004 40328 10080
rect 39988 10964 40328 11040
rect 39988 11924 40328 12000
rect 39988 12884 40328 12960
rect 39988 13844 40328 13920
rect 39988 14804 40328 14880
rect 39988 15764 40328 15840
rect 39988 16724 40328 16800
rect 39988 17684 40328 17760
rect 39988 18644 40328 18720
rect 39988 19604 40328 19680
rect 39988 20564 40328 20640
rect 39988 21524 40328 21600
rect 39988 22484 40328 22560
rect 39988 23444 40328 23520
<< m1 >>
rect 1152 3882 1508 3942
rect 1152 8558 1508 8618
rect 1508 3882 1568 8618
rect 4608 8558 4760 8618
rect 4760 4084 6568 4144
rect 4760 5044 6568 5104
rect 4760 6004 6568 6064
rect 4760 6964 6568 7024
rect 4760 7924 6568 7984
rect 4760 8884 6568 8944
rect 4760 9844 6568 9904
rect 4760 10804 6568 10864
rect 4760 11764 6568 11824
rect 4760 12724 6568 12784
rect 4760 13684 6568 13744
rect 4760 14644 6568 14704
rect 4760 15604 6568 15664
rect 4760 16564 6568 16624
rect 4760 17524 6568 17584
rect 4760 18484 6568 18544
rect 4760 19444 6568 19504
rect 4760 20404 6568 20464
rect 4760 21364 6568 21424
rect 4760 22324 6568 22384
rect 4760 23284 6568 23344
rect 4760 24244 6568 24304
rect 4760 4084 4820 24304
<< m2 >>
rect 4616 3882 4780 3958
rect 4780 1204 6568 1280
rect 4780 2164 6568 2240
rect 4780 3124 6568 3200
rect 4780 1204 4856 3958
use SUNTR_RPPO8 xa1 ../SUN_TR_SKY130NM
transform 1 0 444 0 1 444
box 444 444 5708 4680
use SUNTR_RPPO8 xa2 ../SUN_TR_SKY130NM
transform 1 0 444 0 1 5120
box 444 5120 5708 9356
use CAP_LPF xb1 
transform -1 0 40108 0 1 444
box 40108 444 73788 1404
use CAP_LPF xb2_0 
transform -1 0 40108 0 1 1404
box 40108 1404 73788 2364
use CAP_LPF xb2_1 
transform -1 0 40108 0 1 2364
box 40108 2364 73788 3324
use CAP_LPF xb3_0 
transform -1 0 40108 0 1 3324
box 40108 3324 73788 4284
use CAP_LPF xb3_1 
transform -1 0 40108 0 1 4284
box 40108 4284 73788 5244
use CAP_LPF xb3_10 
transform -1 0 40108 0 1 5244
box 40108 5244 73788 6204
use CAP_LPF xb3_11 
transform -1 0 40108 0 1 6204
box 40108 6204 73788 7164
use CAP_LPF xb3_12 
transform -1 0 40108 0 1 7164
box 40108 7164 73788 8124
use CAP_LPF xb3_13 
transform -1 0 40108 0 1 8124
box 40108 8124 73788 9084
use CAP_LPF xb3_14 
transform -1 0 40108 0 1 9084
box 40108 9084 73788 10044
use CAP_LPF xb3_15 
transform -1 0 40108 0 1 10044
box 40108 10044 73788 11004
use CAP_LPF xb3_16 
transform -1 0 40108 0 1 11004
box 40108 11004 73788 11964
use CAP_LPF xb3_17 
transform -1 0 40108 0 1 11964
box 40108 11964 73788 12924
use CAP_LPF xb3_18 
transform -1 0 40108 0 1 12924
box 40108 12924 73788 13884
use CAP_LPF xb3_19 
transform -1 0 40108 0 1 13884
box 40108 13884 73788 14844
use CAP_LPF xb3_2 
transform -1 0 40108 0 1 14844
box 40108 14844 73788 15804
use CAP_LPF xb3_20 
transform -1 0 40108 0 1 15804
box 40108 15804 73788 16764
use CAP_LPF xb3_21 
transform -1 0 40108 0 1 16764
box 40108 16764 73788 17724
use CAP_LPF xb3_3 
transform -1 0 40108 0 1 17724
box 40108 17724 73788 18684
use CAP_LPF xb3_4 
transform -1 0 40108 0 1 18684
box 40108 18684 73788 19644
use CAP_LPF xb3_5 
transform -1 0 40108 0 1 19644
box 40108 19644 73788 20604
use CAP_LPF xb3_6 
transform -1 0 40108 0 1 20604
box 40108 20604 73788 21564
use CAP_LPF xb3_7 
transform -1 0 40108 0 1 21564
box 40108 21564 73788 22524
use CAP_LPF xb3_8 
transform -1 0 40108 0 1 22524
box 40108 22524 73788 23484
use CAP_LPF xb3_9 
transform -1 0 40108 0 1 23484
box 40108 23484 73788 24444
use cut_M1M4_2x1 xcut0 
transform 1 0 23128 0 1 0
box 23128 0 23328 76
use cut_M1M2_2x1 xcut1 
transform 1 0 1060 0 1 3882
box 1060 3882 1244 3950
use cut_M1M2_2x1 xcut2 
transform 1 0 1060 0 1 8558
box 1060 8558 1244 8626
use cut_M1M2_2x1 xcut3 
transform 1 0 4516 0 1 8558
box 4516 8558 4700 8626
use cut_M2M4_2x1 xcut4 
transform 1 0 6468 0 1 4084
box 6468 4084 6668 4160
use cut_M2M4_2x1 xcut5 
transform 1 0 6468 0 1 5044
box 6468 5044 6668 5120
use cut_M2M4_2x1 xcut6 
transform 1 0 6468 0 1 6004
box 6468 6004 6668 6080
use cut_M2M4_2x1 xcut7 
transform 1 0 6468 0 1 6964
box 6468 6964 6668 7040
use cut_M2M4_2x1 xcut8 
transform 1 0 6468 0 1 7924
box 6468 7924 6668 8000
use cut_M2M4_2x1 xcut9 
transform 1 0 6468 0 1 8884
box 6468 8884 6668 8960
use cut_M2M4_2x1 xcut10 
transform 1 0 6468 0 1 9844
box 6468 9844 6668 9920
use cut_M2M4_2x1 xcut11 
transform 1 0 6468 0 1 10804
box 6468 10804 6668 10880
use cut_M2M4_2x1 xcut12 
transform 1 0 6468 0 1 11764
box 6468 11764 6668 11840
use cut_M2M4_2x1 xcut13 
transform 1 0 6468 0 1 12724
box 6468 12724 6668 12800
use cut_M2M4_2x1 xcut14 
transform 1 0 6468 0 1 13684
box 6468 13684 6668 13760
use cut_M2M4_2x1 xcut15 
transform 1 0 6468 0 1 14644
box 6468 14644 6668 14720
use cut_M2M4_2x1 xcut16 
transform 1 0 6468 0 1 15604
box 6468 15604 6668 15680
use cut_M2M4_2x1 xcut17 
transform 1 0 6468 0 1 16564
box 6468 16564 6668 16640
use cut_M2M4_2x1 xcut18 
transform 1 0 6468 0 1 17524
box 6468 17524 6668 17600
use cut_M2M4_2x1 xcut19 
transform 1 0 6468 0 1 18484
box 6468 18484 6668 18560
use cut_M2M4_2x1 xcut20 
transform 1 0 6468 0 1 19444
box 6468 19444 6668 19520
use cut_M2M4_2x1 xcut21 
transform 1 0 6468 0 1 20404
box 6468 20404 6668 20480
use cut_M2M4_2x1 xcut22 
transform 1 0 6468 0 1 21364
box 6468 21364 6668 21440
use cut_M2M4_2x1 xcut23 
transform 1 0 6468 0 1 22324
box 6468 22324 6668 22400
use cut_M2M4_2x1 xcut24 
transform 1 0 6468 0 1 23284
box 6468 23284 6668 23360
use cut_M2M4_2x1 xcut25 
transform 1 0 6468 0 1 24244
box 6468 24244 6668 24320
use cut_M1M3_2x1 xcut26 
transform 1 0 4516 0 1 3882
box 4516 3882 4716 3958
use cut_M3M4_2x1 xcut27 
transform 1 0 6468 0 1 1204
box 6468 1204 6668 1280
use cut_M3M4_2x1 xcut28 
transform 1 0 6468 0 1 2164
box 6468 2164 6668 2240
use cut_M3M4_2x1 xcut29 
transform 1 0 6468 0 1 3124
box 6468 3124 6668 3200
use cut_M1M4_1x2 xcut30 
transform 1 0 40252 0 1 0
box 40252 0 40328 200
use cut_M1M4_1x2 xcut31 
transform 1 0 40252 0 1 404
box 40252 404 40328 604
use cut_M1M4_1x2 xcut32 
transform 1 0 40252 0 1 1364
box 40252 1364 40328 1564
use cut_M1M4_1x2 xcut33 
transform 1 0 40252 0 1 2324
box 40252 2324 40328 2524
use cut_M1M4_1x2 xcut34 
transform 1 0 40252 0 1 3284
box 40252 3284 40328 3484
use cut_M1M4_1x2 xcut35 
transform 1 0 40252 0 1 4244
box 40252 4244 40328 4444
use cut_M1M4_1x2 xcut36 
transform 1 0 40252 0 1 5204
box 40252 5204 40328 5404
use cut_M1M4_1x2 xcut37 
transform 1 0 40252 0 1 6164
box 40252 6164 40328 6364
use cut_M1M4_1x2 xcut38 
transform 1 0 40252 0 1 7124
box 40252 7124 40328 7324
use cut_M1M4_1x2 xcut39 
transform 1 0 40252 0 1 8084
box 40252 8084 40328 8284
use cut_M1M4_1x2 xcut40 
transform 1 0 40252 0 1 9044
box 40252 9044 40328 9244
use cut_M1M4_1x2 xcut41 
transform 1 0 40252 0 1 10004
box 40252 10004 40328 10204
use cut_M1M4_1x2 xcut42 
transform 1 0 40252 0 1 10964
box 40252 10964 40328 11164
use cut_M1M4_1x2 xcut43 
transform 1 0 40252 0 1 11924
box 40252 11924 40328 12124
use cut_M1M4_1x2 xcut44 
transform 1 0 40252 0 1 12884
box 40252 12884 40328 13084
use cut_M1M4_1x2 xcut45 
transform 1 0 40252 0 1 13844
box 40252 13844 40328 14044
use cut_M1M4_1x2 xcut46 
transform 1 0 40252 0 1 14804
box 40252 14804 40328 15004
use cut_M1M4_1x2 xcut47 
transform 1 0 40252 0 1 15764
box 40252 15764 40328 15964
use cut_M1M4_1x2 xcut48 
transform 1 0 40252 0 1 16724
box 40252 16724 40328 16924
use cut_M1M4_1x2 xcut49 
transform 1 0 40252 0 1 17684
box 40252 17684 40328 17884
use cut_M1M4_1x2 xcut50 
transform 1 0 40252 0 1 18644
box 40252 18644 40328 18844
use cut_M1M4_1x2 xcut51 
transform 1 0 40252 0 1 19604
box 40252 19604 40328 19804
use cut_M1M4_1x2 xcut52 
transform 1 0 40252 0 1 20564
box 40252 20564 40328 20764
use cut_M1M4_1x2 xcut53 
transform 1 0 40252 0 1 21524
box 40252 21524 40328 21724
use cut_M1M4_1x2 xcut54 
transform 1 0 40252 0 1 22484
box 40252 22484 40328 22684
use cut_M1M4_1x2 xcut55 
transform 1 0 40252 0 1 23444
box 40252 23444 40328 23644
<< labels >>
flabel locali s 40252 0 40552 24888 0 FreeSans 400 0 0 0 AVSS
port 2 nsew signal bidirectional
flabel locali s 4516 8558 5092 8778 0 FreeSans 400 0 0 0 VLPFZ
port 1 nsew signal bidirectional
flabel locali s 4516 3882 5092 4102 0 FreeSans 400 0 0 0 VLPF
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 40552 24888
<< end >>
