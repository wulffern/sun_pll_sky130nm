magic
tech sky130B
timestamp 1728046668
<< locali >>
rect 0 12294 20276 12444
rect 0 2624 150 12294
rect 2258 4279 2546 4389
rect 0 2568 230 2624
rect 0 286 150 2568
rect 2258 1941 2546 2051
rect 0 230 230 286
rect 0 150 150 230
rect 20126 150 20276 12294
rect 0 0 20276 150
<< metal1 >>
rect 2380 12122 3284 12152
rect 2380 11672 2410 12122
rect 2380 11642 3284 11672
rect 2380 11192 2410 11642
rect 2380 11162 3284 11192
rect 2380 10712 2410 11162
rect 2380 10682 3284 10712
rect 2380 10232 2410 10682
rect 2380 10202 3284 10232
rect 2380 9752 2410 10202
rect 2380 9722 3284 9752
rect 2380 9272 2410 9722
rect 2380 9242 3284 9272
rect 2380 8792 2410 9242
rect 2380 8762 3284 8792
rect 2380 8312 2410 8762
rect 2380 8282 3284 8312
rect 2380 7832 2410 8282
rect 2380 7802 3284 7832
rect 2380 7352 2410 7802
rect 2380 7322 3284 7352
rect 2380 6872 2410 7322
rect 2380 6842 3284 6872
rect 2380 6392 2410 6842
rect 2380 6362 3284 6392
rect 2380 5912 2410 6362
rect 2380 5882 3284 5912
rect 2380 5432 2410 5882
rect 2380 5402 3284 5432
rect 2380 4952 2410 5402
rect 2380 4922 3284 4952
rect 2380 4472 2410 4922
rect 2380 4442 3284 4472
rect 2380 4309 2410 4442
rect 576 4279 784 4309
rect 2304 4279 2410 4309
rect 754 1971 784 4279
rect 2380 3992 2410 4279
rect 2380 3962 3284 3992
rect 2380 3512 2410 3962
rect 2380 3482 3284 3512
rect 2380 3032 2410 3482
rect 2380 3002 3284 3032
rect 2380 2552 2410 3002
rect 2380 2522 3284 2552
rect 2380 2072 2410 2522
rect 2380 2042 3284 2072
rect 576 1941 784 1971
<< metal2 >>
rect 2308 1941 2428 1979
rect 2390 1600 2428 1941
rect 2390 1562 3284 1600
rect 2390 1120 2428 1562
rect 2390 1082 3284 1120
rect 2390 640 2428 1082
rect 2390 602 3284 640
<< metal3 >>
rect 19994 11722 20164 11760
rect 19994 11242 20164 11280
rect 19994 10762 20164 10800
rect 19994 10282 20164 10320
rect 19994 9802 20164 9840
rect 19994 9322 20164 9360
rect 19994 8842 20164 8880
rect 19994 8362 20164 8400
rect 19994 7882 20164 7920
rect 19994 7402 20164 7440
rect 19994 6922 20164 6960
rect 19994 6442 20164 6480
rect 19994 5962 20164 6000
rect 19994 5482 20164 5520
rect 19994 5002 20164 5040
rect 19994 4522 20164 4560
rect 19994 4042 20164 4080
rect 19994 3562 20164 3600
rect 19994 3082 20164 3120
rect 19994 2602 20164 2640
rect 19994 2122 20164 2160
rect 19994 1642 20164 1680
rect 19994 1162 20164 1200
rect 19994 682 20164 720
rect 11560 0 11668 242
rect 19994 202 20164 240
use SUNTR_RPPO8  xa1 ../SUN_TR_SKY130NM
timestamp 1728046668
transform 1 0 222 0 1 222
box 0 0 2632 2118
use SUNTR_RPPO8  xa2
timestamp 1728046668
transform 1 0 222 0 1 2560
box 0 0 2632 2118
use CAP_LPF  xb1
timestamp 1720908000
transform -1 0 20054 0 1 222
box 60 -20 16820 420
use CAP_LPF  xb2_0
timestamp 1720908000
transform -1 0 20054 0 1 702
box 60 -20 16820 420
use CAP_LPF  xb2_1
timestamp 1720908000
transform -1 0 20054 0 1 1182
box 60 -20 16820 420
use CAP_LPF  xb3_0
timestamp 1720908000
transform -1 0 20054 0 1 1662
box 60 -20 16820 420
use CAP_LPF  xb3_1
timestamp 1720908000
transform -1 0 20054 0 1 2142
box 60 -20 16820 420
use CAP_LPF  xb3_2
timestamp 1720908000
transform -1 0 20054 0 1 7422
box 60 -20 16820 420
use CAP_LPF  xb3_3
timestamp 1720908000
transform -1 0 20054 0 1 8862
box 60 -20 16820 420
use CAP_LPF  xb3_4
timestamp 1720908000
transform -1 0 20054 0 1 9342
box 60 -20 16820 420
use CAP_LPF  xb3_5
timestamp 1720908000
transform -1 0 20054 0 1 9822
box 60 -20 16820 420
use CAP_LPF  xb3_6
timestamp 1720908000
transform -1 0 20054 0 1 10302
box 60 -20 16820 420
use CAP_LPF  xb3_7
timestamp 1720908000
transform -1 0 20054 0 1 10782
box 60 -20 16820 420
use CAP_LPF  xb3_8
timestamp 1720908000
transform -1 0 20054 0 1 11262
box 60 -20 16820 420
use CAP_LPF  xb3_9
timestamp 1720908000
transform -1 0 20054 0 1 11742
box 60 -20 16820 420
use CAP_LPF  xb3_10
timestamp 1720908000
transform -1 0 20054 0 1 2622
box 60 -20 16820 420
use CAP_LPF  xb3_11
timestamp 1720908000
transform -1 0 20054 0 1 3102
box 60 -20 16820 420
use CAP_LPF  xb3_12
timestamp 1720908000
transform -1 0 20054 0 1 3582
box 60 -20 16820 420
use CAP_LPF  xb3_13
timestamp 1720908000
transform -1 0 20054 0 1 4062
box 60 -20 16820 420
use CAP_LPF  xb3_14
timestamp 1720908000
transform -1 0 20054 0 1 4542
box 60 -20 16820 420
use CAP_LPF  xb3_15
timestamp 1720908000
transform -1 0 20054 0 1 5022
box 60 -20 16820 420
use CAP_LPF  xb3_16
timestamp 1720908000
transform -1 0 20054 0 1 5502
box 60 -20 16820 420
use CAP_LPF  xb3_17
timestamp 1720908000
transform -1 0 20054 0 1 5982
box 60 -20 16820 420
use CAP_LPF  xb3_18
timestamp 1720908000
transform -1 0 20054 0 1 6462
box 60 -20 16820 420
use CAP_LPF  xb3_19
timestamp 1720908000
transform -1 0 20054 0 1 6942
box 60 -20 16820 420
use CAP_LPF  xb3_20
timestamp 1720908000
transform -1 0 20054 0 1 7902
box 60 -20 16820 420
use CAP_LPF  xb3_21
timestamp 1720908000
transform -1 0 20054 0 1 8382
box 60 -20 16820 420
use cut_M1M4_2x1  xcut0
timestamp 1720908000
transform 1 0 11564 0 1 0
box 0 0 100 38
use cut_M1M2_2x1  xcut1
timestamp 1720908000
transform 1 0 530 0 1 1941
box 0 0 92 34
use cut_M1M2_2x1  xcut2
timestamp 1720908000
transform 1 0 530 0 1 4279
box 0 0 92 34
use cut_M1M2_2x1  xcut3
timestamp 1720908000
transform 1 0 2258 0 1 4279
box 0 0 92 34
use cut_M2M4_2x1  xcut4
timestamp 1720908000
transform 1 0 3234 0 1 2042
box 0 0 100 38
use cut_M2M4_2x1  xcut5
timestamp 1720908000
transform 1 0 3234 0 1 2522
box 0 0 100 38
use cut_M2M4_2x1  xcut6
timestamp 1720908000
transform 1 0 3234 0 1 3002
box 0 0 100 38
use cut_M2M4_2x1  xcut7
timestamp 1720908000
transform 1 0 3234 0 1 3482
box 0 0 100 38
use cut_M2M4_2x1  xcut8
timestamp 1720908000
transform 1 0 3234 0 1 3962
box 0 0 100 38
use cut_M2M4_2x1  xcut9
timestamp 1720908000
transform 1 0 3234 0 1 4442
box 0 0 100 38
use cut_M2M4_2x1  xcut10
timestamp 1720908000
transform 1 0 3234 0 1 4922
box 0 0 100 38
use cut_M2M4_2x1  xcut11
timestamp 1720908000
transform 1 0 3234 0 1 5402
box 0 0 100 38
use cut_M2M4_2x1  xcut12
timestamp 1720908000
transform 1 0 3234 0 1 5882
box 0 0 100 38
use cut_M2M4_2x1  xcut13
timestamp 1720908000
transform 1 0 3234 0 1 6362
box 0 0 100 38
use cut_M2M4_2x1  xcut14
timestamp 1720908000
transform 1 0 3234 0 1 6842
box 0 0 100 38
use cut_M2M4_2x1  xcut15
timestamp 1720908000
transform 1 0 3234 0 1 7322
box 0 0 100 38
use cut_M2M4_2x1  xcut16
timestamp 1720908000
transform 1 0 3234 0 1 7802
box 0 0 100 38
use cut_M2M4_2x1  xcut17
timestamp 1720908000
transform 1 0 3234 0 1 8282
box 0 0 100 38
use cut_M2M4_2x1  xcut18
timestamp 1720908000
transform 1 0 3234 0 1 8762
box 0 0 100 38
use cut_M2M4_2x1  xcut19
timestamp 1720908000
transform 1 0 3234 0 1 9242
box 0 0 100 38
use cut_M2M4_2x1  xcut20
timestamp 1720908000
transform 1 0 3234 0 1 9722
box 0 0 100 38
use cut_M2M4_2x1  xcut21
timestamp 1720908000
transform 1 0 3234 0 1 10202
box 0 0 100 38
use cut_M2M4_2x1  xcut22
timestamp 1720908000
transform 1 0 3234 0 1 10682
box 0 0 100 38
use cut_M2M4_2x1  xcut23
timestamp 1720908000
transform 1 0 3234 0 1 11162
box 0 0 100 38
use cut_M2M4_2x1  xcut24
timestamp 1720908000
transform 1 0 3234 0 1 11642
box 0 0 100 38
use cut_M2M4_2x1  xcut25
timestamp 1720908000
transform 1 0 3234 0 1 12122
box 0 0 100 38
use cut_M1M3_2x1  xcut26
timestamp 1720908000
transform 1 0 2258 0 1 1941
box 0 0 100 38
use cut_M3M4_2x1  xcut27
timestamp 1720908000
transform 1 0 3234 0 1 602
box 0 0 100 38
use cut_M3M4_2x1  xcut28
timestamp 1720908000
transform 1 0 3234 0 1 1082
box 0 0 100 38
use cut_M3M4_2x1  xcut29
timestamp 1720908000
transform 1 0 3234 0 1 1562
box 0 0 100 38
use cut_M1M4_1x2  xcut30
timestamp 1720908000
transform 1 0 20126 0 1 0
box 0 0 38 100
use cut_M1M4_1x2  xcut31
timestamp 1720908000
transform 1 0 20126 0 1 202
box 0 0 38 100
use cut_M1M4_1x2  xcut32
timestamp 1720908000
transform 1 0 20126 0 1 682
box 0 0 38 100
use cut_M1M4_1x2  xcut33
timestamp 1720908000
transform 1 0 20126 0 1 1162
box 0 0 38 100
use cut_M1M4_1x2  xcut34
timestamp 1720908000
transform 1 0 20126 0 1 1642
box 0 0 38 100
use cut_M1M4_1x2  xcut35
timestamp 1720908000
transform 1 0 20126 0 1 2122
box 0 0 38 100
use cut_M1M4_1x2  xcut36
timestamp 1720908000
transform 1 0 20126 0 1 2602
box 0 0 38 100
use cut_M1M4_1x2  xcut37
timestamp 1720908000
transform 1 0 20126 0 1 3082
box 0 0 38 100
use cut_M1M4_1x2  xcut38
timestamp 1720908000
transform 1 0 20126 0 1 3562
box 0 0 38 100
use cut_M1M4_1x2  xcut39
timestamp 1720908000
transform 1 0 20126 0 1 4042
box 0 0 38 100
use cut_M1M4_1x2  xcut40
timestamp 1720908000
transform 1 0 20126 0 1 4522
box 0 0 38 100
use cut_M1M4_1x2  xcut41
timestamp 1720908000
transform 1 0 20126 0 1 5002
box 0 0 38 100
use cut_M1M4_1x2  xcut42
timestamp 1720908000
transform 1 0 20126 0 1 5482
box 0 0 38 100
use cut_M1M4_1x2  xcut43
timestamp 1720908000
transform 1 0 20126 0 1 5962
box 0 0 38 100
use cut_M1M4_1x2  xcut44
timestamp 1720908000
transform 1 0 20126 0 1 6442
box 0 0 38 100
use cut_M1M4_1x2  xcut45
timestamp 1720908000
transform 1 0 20126 0 1 6922
box 0 0 38 100
use cut_M1M4_1x2  xcut46
timestamp 1720908000
transform 1 0 20126 0 1 7402
box 0 0 38 100
use cut_M1M4_1x2  xcut47
timestamp 1720908000
transform 1 0 20126 0 1 7882
box 0 0 38 100
use cut_M1M4_1x2  xcut48
timestamp 1720908000
transform 1 0 20126 0 1 8362
box 0 0 38 100
use cut_M1M4_1x2  xcut49
timestamp 1720908000
transform 1 0 20126 0 1 8842
box 0 0 38 100
use cut_M1M4_1x2  xcut50
timestamp 1720908000
transform 1 0 20126 0 1 9322
box 0 0 38 100
use cut_M1M4_1x2  xcut51
timestamp 1720908000
transform 1 0 20126 0 1 9802
box 0 0 38 100
use cut_M1M4_1x2  xcut52
timestamp 1720908000
transform 1 0 20126 0 1 10282
box 0 0 38 100
use cut_M1M4_1x2  xcut53
timestamp 1720908000
transform 1 0 20126 0 1 10762
box 0 0 38 100
use cut_M1M4_1x2  xcut54
timestamp 1720908000
transform 1 0 20126 0 1 11242
box 0 0 38 100
use cut_M1M4_1x2  xcut55
timestamp 1720908000
transform 1 0 20126 0 1 11722
box 0 0 38 100
<< labels >>
flabel locali s 20126 0 20276 12444 0 FreeSans 400 0 0 0 AVSS
port 2 nsew signal bidirectional
flabel locali s 2258 4279 2546 4389 0 FreeSans 400 0 0 0 VLPFZ
port 1 nsew signal bidirectional
flabel locali s 2258 1941 2546 2051 0 FreeSans 400 0 0 0 VLPF
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 20276 12444
<< end >>
