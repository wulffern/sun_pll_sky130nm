* NGSPICE file created from SUN_PLL.ext - technology: sky130B

.subckt SUN_PLL PWRUP_1V8 CK_REF CK IBPSR_1U AVSS AVDD
X0 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R0 AVSS m3_37748_115804# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X1 xaa1.xa2.M8.D IBPSR_1U xaa1.xa2.M7.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R1 m3_4628_94524# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X2 xaa4.xa1.M6.D IBPSR_1U xaa4.xa1.M5.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X3 xaa6.xf.XA6.MN0.G xaa6.xf.XA5.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R2 AVSS m3_37748_107164# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X4 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=73.5 pd=387 as=0.616 ps=3.3 w=1.08 l=0.18
X5 xaa6.xf.XA7.MN1.G PWRUP_1V8 xaa6.xf.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X6 xaa0.xa3.MP0.D xaa0.xa1.MN2.S AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X7 AVDD PWRUP_1V8 xaa6.xd.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X8 xaa6.xe.XA7.MP1.G xaa6.xe.XA7.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X9 xaa5.xb2_1.MN0.D xaa5.xb2_0.MN0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X10 xaa6.xd.XA5.MN0.G xaa6.xd.XA7.MP1.G xaa6.xd.XA3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X11 xaa6.xf.XA5.MN0.G xaa6.xf.XA7.MP1.G xaa6.xf.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X12 xaa3.xa5a.MN0.D xaa3.xa4.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X13 AVDD xaa4.xa2.M0.D xaa4.xa4.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X14 xaa4.xa1.M8.D IBPSR_1U xaa4.xa1.M7.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R3 AVSS m3_37748_78364# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X15 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MN1.G xaa6.xe.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R4 AVSS m3_37748_102364# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X16 xaa5.xb3.MP1.D xaa5.xb3.MP1.D xaa5.xb3.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=1.23 pd=6.6 as=0.616 ps=3.3 w=1.08 l=0.18
R5 AVSS m3_37748_99484# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X17 xaa3.xa4.MN0.D xaa3.xa3a.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R6 m3_4628_81084# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R7 m3_4628_116604# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X18 xaa6.xe.XA3.MP0.D xaa6.xe.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X19 xaa6.xd.XA4.MP0.D xaa6.xd.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X20 a_2084_70022# xaa1.xa3.D AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X21 xaa5.xb2_2.MN0.D xaa5.xb2_1.MN0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X22 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X23 xaa6.xe.XA6.MP0.D xaa6.xe.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X24 xaa5.xb1.MN1.G xaa5.xa3.xb1_0.G xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R8 AVSS m3_37748_73564# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X25 xaa6.xc.XA7.MP1.G xaa6.xc.XA7.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X26 xaa1.xa2.M7.D IBPSR_1U xaa1.xa2.M6.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X27 xaa1.xa1.M5.D IBPSR_1U xaa1.xa1.M4.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R9 m3_4628_89724# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X28 xaa1.xb2.M0.D xaa1.xa1.M8.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
R10 AVSS m3_37748_94684# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R11 m3_4628_111804# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X29 a_356_74698# a_n76_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X30 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MP1.G xaa6.xc.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X31 xaa1.xa2.M5.D IBPSR_1U xaa1.xa2.M4.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X32 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R12 m3_4628_103164# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X33 xaa6.xc.XA3.MN0.D xaa6.xc.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X34 xaa5.xa3.xb2_0.D xaa5.xa3.xb2_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X35 xaa1.xa1.M3.D IBPSR_1U xaa1.xa1.M2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R13 AVSS li_6204_57236# sky130_fd_pr__res_generic_l1 w=0.44 l=0.36
X36 a_n508_70022# xbb0.xa1.XA1.N AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X37 xaa3.xa2.MN0.D xaa3.xa1capd.B AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X38 a_2084_74698# a_1652_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X39 xaa6.xc.XA6.MN0.D xaa6.xc.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R14 m3_4628_84924# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X40 xaa6.xf.XA7.MP1.G xaa6.xf.XA7.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X41 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=61.6 pd=330 as=0.616 ps=3.3 w=1.08 l=0.18
X42 xaa4.xa1.M5.D IBPSR_1U xaa4.xa1.M4.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R15 m3_4628_76284# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X43 xaa6.xd.XA7.MN2.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X44 xaa6.xd.XA5.MN0.G xaa6.xd.XA7.MN1.G xaa6.xd.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X45 xaa5.xb2_1.MN0.D xaa5.xb2_0.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X46 xaa3.xa3a.MN0.D xaa3.xa2.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R16 xaa4.xa2.M0.G m3_22620_60292# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X47 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MN1.G xaa6.xf.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R17 AVSS m3_37748_86044# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X48 xaa4.xa4.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X49 xaa4.xa1.M3.D IBPSR_1U xaa4.xa1.M2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X50 xaa1.xa4.M0.G xaa3.xa7.MN0.D xaa3.xa8.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X51 xaa6.xf.XA3.MP0.D xaa6.xf.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R18 AVSS m3_37748_110044# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X52 IBPSR_1U IBPSR_1U xbb1.xa3.M7.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X53 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R19 AVSS m3_37748_89884# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R20 m3_4628_71484# xaa1.xa3.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X54 xaa6.xf.XA6.MP0.D xaa6.xf.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X55 xaa5.xa3.xc1a.D xaa5.xa3.xb2_0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X56 xaa6.xd.XA4.MN0.D xaa6.xd.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X57 xaa5.xb2_2.MN0.D xaa5.xb2_1.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R21 AVSS m3_37748_113884# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X58 xaa6.xg.XA1.MN0.D CK AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X59 xaa3.xa7.MN0.D xaa3.xa6.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X60 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X61 CK xaa5.xa3.xb2_0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X62 xaa0.xa1.MN0.D xaa0.xa1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X63 xbb1.xa3.M6.D IBPSR_1U xbb1.xa3.M5.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X64 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X65 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X66 xaa5.xb1.MN1.G xaa5.xa3.xb1_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R22 AVSS m3_37748_81244# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R23 m3_13044_61524# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X67 AVDD PWRUP_1V8 xaa6.xg.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X68 xaa6.xc.XA7.MN1.G xaa6.xc.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X69 xaa6.xe.XA6.MN0.G xaa6.xe.XA5.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X70 xaa6.xg.XA5.MN0.G xaa6.xg.XA7.MP1.G xaa6.xg.XA3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R24 m3_4628_97404# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X71 xaa6.xe.XA7.MN1.G PWRUP_1V8 xaa6.xe.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X72 xaa1.xa4.M0.D xaa1.xa4.M0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X73 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X74 xaa3.xa1b.MN0.D PWRUP_1V8 AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X75 xaa1.xa4.M0.G xaa3.xa1b.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X76 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X77 xaa1.xa2.M0.D IBPSR_1U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X78 xaa6.xe.XA5.MN0.G xaa6.xe.XA7.MP1.G xaa6.xe.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X79 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X80 a_1220_70022# a_1652_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R25 m3_13044_55188# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X81 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MN1.G xaa6.xg.XA7.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X82 xaa6.xg.XA4.MP0.D xaa6.xg.XA4.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R26 m3_13044_58356# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R27 m3_4628_92604# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R28 m3_4628_114684# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X83 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MP1.G xaa6.xc.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R29 xaa4.xa2.M0.G m3_22620_57124# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X84 xaa6.xf.XA7.MP1.G xaa6.xf.XA7.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R30 AVSS m3_37748_105244# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X85 xaa1.xa2.M2.D IBPSR_1U xaa1.xa2.M1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X86 xaa4.xa1.M0.D IBPSR_1U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X87 xaa6.xg.XA7.MN0.D xaa6.xg.XA7.MN0.G xaa6.xg.XA7.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X88 xaa0.xa1.MP1.D xaa0.xa1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X89 xaa6.xc.XA7.MN0.D xaa0.xa5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X90 xaa4.xa2.M0.D xaa4.xa2.M0.G xaa4.xa1.M8.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X91 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MP1.G xaa6.xf.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R31 AVSS m3_37748_76444# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X92 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X93 xaa5.xb1.MN1.D PWRUP_1V8 xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X94 xaa6.xf.XA3.MN0.D xaa6.xf.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X95 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X96 AVDD PWRUP_1V8 xaa6.xe.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R32 AVSS m3_37748_100444# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X97 xbb1.xa3.M3.D IBPSR_1U xbb1.xa3.M2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R33 AVSS m3_37748_97564# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X98 xaa6.xe.XA5.MN0.G xaa6.xe.XA7.MP1.G xaa6.xe.XA3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X99 xaa5.xb2_3.MN0.D xaa5.xb2_2.MN0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X100 xaa6.xf.XA6.MN0.D xaa6.xf.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X101 xaa6.xd.XA7.MN1.G xaa6.xd.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R34 m3_4628_106044# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X102 xbb1.xa3.M1.D IBPSR_1U xbb1.xa3.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X103 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R35 AVSS m3_37748_71644# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X104 xaa6.xe.XA4.MP0.D xaa6.xe.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X105 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X106 xaa5.xb2_4.MN0.D xaa5.xb2_3.MN0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R36 m3_4628_87804# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R37 m3_4628_109884# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X107 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X108 xaa3.xa5a.MN0.D xaa3.xa4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X109 xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
R38 AVSS m3_37748_92764# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X110 xaa6.xc.XA7.MN2.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R39 m3_4628_79164# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X111 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X112 xaa6.xc.XA5.MN0.G xaa6.xc.XA7.MN1.G xaa6.xc.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X113 xaa5.xa3.xb2_0.D xaa5.xa3.xb2_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X114 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R40 m3_4628_101244# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X115 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MP1.G xaa6.xd.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X116 xaa3.xa4.MN0.D xaa3.xa3a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X117 xaa6.xd.XA7.MN0.D xaa6.xc.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X118 xaa6.xc.XA4.MN0.D xaa6.xc.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X119 xaa5.xa4.MN0.D xaa5.xa3.xb1_0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X120 xaa1.xa1.M7.D IBPSR_1U xaa1.xa1.M6.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R41 m3_4628_74364# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X121 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R42 AVSS m3_37748_116764# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X122 AVDD PWRUP_1V8 xaa6.xf.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R43 m3_4628_95484# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R44 AVSS m3_37748_84124# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X123 xaa6.xf.XA5.MN0.G xaa6.xf.XA7.MP1.G xaa6.xf.XA3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X124 xaa5.xb1.MN0.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X125 IBPSR_1U xaa3.xa1b.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X126 a_356_70022# a_n76_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X127 xaa5.xb2_3.MN0.D xaa5.xb2_2.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R45 AVSS m3_37748_87964# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X128 xaa6.xd.XA1.MN0.D xaa6.xd.XA1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X129 xaa4.xa1.M7.D IBPSR_1U xaa4.xa1.M6.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R46 AVSS m3_37748_111964# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X130 xaa6.xf.XA4.MP0.D xaa6.xf.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X131 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X132 a_356_74698# a_788_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R47 m3_4628_90684# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X133 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X134 a_2084_70022# a_1652_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R48 m3_4628_117564# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X135 xaa6.xe.XA7.MP1.G xaa6.xe.XA7.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X136 AVDD xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X137 xaa5.xb2_4.MN0.D xaa5.xb2_3.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R49 m3_13044_54132# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R50 AVSS m3_37748_108124# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X138 xaa4.xa4.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X139 xaa3.xa9.MN0.D xaa1.xa4.M0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X140 AVSS xaa3.xa7.MN0.D xaa1.xa4.M0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R51 m3_13044_57300# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R52 m3_4628_69564# xaa1.xa3.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X141 xaa5.xa3.xb1_0.D xaa5.xa3.xb2_0.D xaa5.xa3.xc1a.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X142 AVDD xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X143 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MP1.G xaa6.xe.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X144 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MN1.G xaa6.xd.XA7.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X145 xaa6.xf.XA1.MN0.G xaa6.xg.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X146 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X147 xaa6.xg.XA3.MN1.G CK AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X148 xaa6.xe.XA3.MN0.D xaa6.xe.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X149 xaa6.xg.XA5.MN0.D xaa6.xg.XA5.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R53 AVSS m3_37748_79324# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X150 xaa0.xa5.MN0.D xaa0.xa1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X151 xaa0.xa5.MN2.G xaa6.xc.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X152 xaa6.xg.XA3.MN1.G PWRUP_1V8 xaa6.xg.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X153 a_n508_74698# a_n76_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R54 m3_4628_112764# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X154 xaa6.xc.XA6.MN0.G xaa6.xc.XA5.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X155 xaa0.xa1.MN2.D CK_REF xaa0.xa1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X156 xaa6.xe.XA6.MN0.D xaa6.xe.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X157 xaa6.xd.XA7.MN0.D xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R55 AVSS m3_37748_103324# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X158 AVDD PWRUP_1V8 xaa6.xc.XA7.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R56 m3_4628_82044# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X159 xaa6.xg.XA5.MN0.G xaa6.xg.XA7.MP1.G xaa6.xg.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X160 xaa1.xa1.M2.D IBPSR_1U xaa1.xa1.M1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X161 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X162 AVSS xaa0.xa3.MN1.G xaa0.xa1.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X163 xaa6.xf.XA7.MN2.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X164 xaa6.xc.XA5.MN0.G xaa6.xc.XA7.MN1.G xaa6.xc.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R57 m3_4628_85884# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X165 xaa6.xf.XA5.MN0.G xaa6.xf.XA7.MN1.G xaa6.xf.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X166 xaa3.xa1b.MN0.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R58 AVSS m3_37748_74524# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X167 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MP1.G xaa6.xg.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X168 xbb1.xa3.M5.D IBPSR_1U xbb1.xa3.M4.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R59 AVSS m3_37748_95644# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X169 xaa4.xa1.M2.D IBPSR_1U xaa4.xa1.M1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X170 xaa6.xg.XA7.MN0.D xaa6.xg.XA7.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X171 xaa6.xf.XA4.MN0.D xaa6.xf.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R60 m3_4628_104124# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X172 xaa0.xa5.MP1.D xaa0.xa1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X173 xbb1.xa3.M7.D IBPSR_1U xbb1.xa3.M6.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X174 xaa0.xa1.MN0.D CK_REF xaa0.xa1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X175 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X176 xaa6.xe.XA7.MN1.G xaa6.xe.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X177 xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R61 m3_4628_107964# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X178 xaa3.xa1capd.B xaa3.xa1b.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X179 xaa4.xa2.M0.G xaa5.xb1.MN1.G xaa5.xb1.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X180 xaa0.xa1.MN0.G xaa0.xa3.MN1.G xaa0.xa3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R62 AVSS m3_37748_90844# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R63 m3_4628_77244# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X181 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X182 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X183 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X184 xaa6.xd.XA6.MN0.G xaa6.xd.XA5.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R64 m3_4628_98364# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X185 xaa5.xa3.xb1_0.D xaa5.xa3.xb1_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X186 xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R65 AVSS m3_37748_87004# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X187 AVDD PWRUP_1V8 xaa6.xd.XA7.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R66 AVSS m3_37748_69724# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X188 AVDD xaa4.xa2.M0.D xaa4.xa4.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X189 CK xaa5.xa3.xb2_0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R67 AVSS m3_37748_111004# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X190 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MP1.G xaa6.xe.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X191 xaa6.xd.XA5.MN0.G xaa6.xd.XA7.MN1.G xaa6.xd.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X192 xaa6.xc.XA1.MN0.D xaa6.xc.XA1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R68 m3_4628_72444# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R69 m3_13044_60468# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R70 AVSS m3_37748_114844# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R71 m3_4628_93564# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X193 xaa6.xe.XA7.MN0.D xaa6.xd.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R72 AVSS m3_37748_82204# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X194 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X195 a_1220_74698# a_788_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X196 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MN1.G xaa6.xc.XA7.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X197 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R73 xaa4.xa2.M0.G m3_22620_56068# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X198 xaa6.xf.XA7.MN1.G xaa6.xf.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R74 xaa4.xa2.M0.G m3_22620_59236# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X199 xbb1.xa3.M2.D IBPSR_1U xbb1.xa3.M1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X200 xaa1.xb1.M0.D xaa1.xa1.M8.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X201 xaa6.xc.XA7.MN0.D xaa0.xa5.MN2.G xaa6.xc.XA7.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R75 m3_4628_115644# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X202 xaa4.xa4.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X203 xaa5.xb1.MN1.D xaa5.xb1.MN1.G xaa5.xb1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R76 AVSS m3_37748_106204# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X204 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X205 xbb1.xa3.M0.D IBPSR_1U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X206 xaa6.xe.XA7.MN2.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X207 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X208 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X209 xaa1.xa1.M0.D IBPSR_1U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X210 xaa6.xe.XA5.MN0.G xaa6.xe.XA7.MN1.G xaa6.xe.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X211 xaa6.xd.XA6.MN0.G xaa6.xd.XA5.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X212 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R77 m3_4628_88764# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X213 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MP1.G xaa6.xf.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X214 xaa6.xd.XA7.MN1.G PWRUP_1V8 xaa6.xd.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X215 xaa6.xg.XA7.MP1.G xaa6.xg.XA3.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R78 AVSS m3_37748_77404# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X216 AVSS xaa0.xa1.MN0.D xaa0.xa1.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R79 m3_4628_110844# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X217 xaa3.xa6.MN0.D xaa3.xa5a.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X218 xaa6.xc.XA7.MP1.G xaa6.xc.XA7.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R80 AVSS m3_37748_101404# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X219 xaa6.xd.XA5.MN0.G xaa6.xd.XA7.MP1.G xaa6.xd.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X220 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
R81 AVSS m3_37748_98524# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R82 m3_4628_80124# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X221 xaa6.xf.XA7.MN0.D xaa6.xe.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R83 xaa4.xa2.M0.G m3_22620_53956# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X222 xaa6.xe.XA4.MN0.D xaa6.xe.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X223 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MP1.G xaa6.xg.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X224 a_356_70022# a_788_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X225 AVSS xaa0.xa5.MN0.D xaa0.xa5.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X226 xaa6.xg.XA3.MN0.D xaa6.xg.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R84 m3_4628_107004# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X227 xaa3.xa9.MN0.D xaa1.xa4.M0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R85 m3_4628_83964# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X228 xaa0.xa2a.MN0.G xaa0.xa1.MN2.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X229 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MN1.G xaa6.xc.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X230 xaa6.xf.XA1.MN0.G xaa6.xg.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R86 AVSS m3_37748_72604# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X231 xaa6.xc.XA3.MP0.D xaa6.xc.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X232 xaa5.xa3.xc2a.D xaa5.xa3.xb1_0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X233 xaa6.xg.XA6.MN0.D xaa6.xg.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X234 xaa6.xg.XA5.MN0.D xaa6.xg.XA5.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X235 xaa1.xb2.M7.D xaa1.xa1.M8.D xaa1.xb2.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X236 xaa0.xa5.MN2.D xaa0.xa5.MN2.G xaa0.xa3.MN1.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X237 AVDD PWRUP_1V8 xaa6.xg.XA3.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R87 AVSS m3_37748_93724# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X238 xaa6.xc.XA6.MP0.D xaa6.xc.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X239 xaa1.xa2.M6.D IBPSR_1U xaa1.xa2.M5.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R88 AVSS m3_37748_85084# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X240 xaa6.xg.XA5.MN0.G xaa6.xg.XA4.MP1.G xaa6.xg.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R89 m3_4628_102204# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X241 xaa6.xf.XA1.MN0.D xaa6.xf.XA1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X242 xaa0.xa1.MN2.S xaa0.xa1.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X243 xaa1.xa1.M4.D IBPSR_1U xaa1.xa1.M3.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R90 AVSS li_6204_59524# sky130_fd_pr__res_generic_l1 w=0.44 l=0.36
X244 a_n508_70022# a_n76_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X245 xaa1.xa2.M4.D IBPSR_1U xaa1.xa2.M3.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X246 xaa0.xa3.MN1.G xaa0.xa5.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X247 a_2084_74698# xaa1.xa4.M0.D AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X248 AVDD xaa4.xa2.M0.D xaa4.xa4.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R91 m3_4628_75324# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X249 xaa0.xa2a.MN0.G xaa0.xa1.MN2.S AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X250 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
R92 AVSS m3_37748_80284# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R93 li_4836_58996# xaa3.xa3a.MN0.D sky130_fd_pr__res_generic_l1 w=0.44 l=0.36
R94 AVSS m3_37748_117724# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X251 xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R95 m3_4628_96444# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X252 xaa6.xd.XA7.MP1.G xaa6.xd.XA7.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X253 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MN1.G xaa6.xf.XA7.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X254 xaa0.xa5.MN0.D xaa0.xa5.MN2.G xaa0.xa5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R96 xaa4.xa2.M0.G m3_22620_58180# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X255 AVDD xaa4.xa2.M0.D xaa4.xa4.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X256 xaa4.xa1.M4.D IBPSR_1U xaa4.xa1.M3.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R97 AVSS m3_37748_109084# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X257 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X258 xaa4.xa1.M8.D xaa1.xa3.D xaa4.xa4.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X259 xaa6.xe.XA6.MN0.G xaa6.xe.XA5.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R98 AVSS m3_37748_88924# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X260 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MN1.G xaa6.xd.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X261 xaa5.xa3.xb1_0.G xaa5.xa3.xb2_0.G xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R99 m3_4628_70524# xaa1.xa3.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X262 xaa6.xf.XA7.MN0.D xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X263 AVDD PWRUP_1V8 xaa6.xe.XA7.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X264 xaa6.xd.XA3.MP0.D xaa6.xd.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X265 xaa3.xa1capd.B xaa3.xa1b.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X266 xaa5.xb2_0.MN0.D xaa5.xb1.MN1.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R100 AVSS m3_37748_112924# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R101 m3_4628_91644# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X267 a_n508_74698# xbb0.xa1.XA1.N AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R102 m3_13044_53076# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X268 xaa6.xe.XA5.MN0.G xaa6.xe.XA7.MN1.G xaa6.xe.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R103 m3_13044_56244# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X269 xaa6.xd.XA6.MP0.D xaa6.xd.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X270 xaa5.xa3.xb2_0.G xaa5.xb2_4.MN0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R104 AVSS m3_37748_104284# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R105 m3_13044_59412# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X271 xaa5.xa3.xb1_0.D xaa5.xa3.xb1_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R106 xaa4.xa2.M0.G m3_22620_55012# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X272 xaa3.xa2.MN0.D xaa3.xa1capd.B AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X273 xaa0.xa5.MN2.G xaa6.xc.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X274 AVSS xaa1.xa4.M0.G xaa1.xa4.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X275 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X276 xaa6.xc.XA6.MN0.G xaa6.xc.XA5.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X277 xaa1.xa2.M1.D IBPSR_1U xaa1.xa2.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R107 AVSS m3_37748_75484# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X278 xbb1.xa3.M4.D IBPSR_1U xbb1.xa3.M3.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X279 xaa6.xc.XA7.MN1.G PWRUP_1V8 xaa6.xc.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X280 xaa1.xa1.M8.D xaa1.xa1.M8.D xaa1.xb1.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X281 xaa3.xa3a.MN0.D xaa3.xa2.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R108 m3_4628_113724# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X282 xaa6.xc.XA5.MN0.G xaa6.xc.XA7.MP1.G xaa6.xc.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X283 xaa1.xa2.M3.D IBPSR_1U xaa1.xa2.M2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R109 m3_4628_105084# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R110 m3_4628_83004# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X284 xaa4.xa4.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X285 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R111 AVSS m3_37748_70684# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X286 xaa1.xa1.M1.D IBPSR_1U xaa1.xa1.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X287 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X288 xaa6.xd.XA7.MP1.G xaa6.xd.XA7.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X289 AVDD xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X290 xaa4.xa1.M8.D xaa4.xa2.M0.G xaa4.xa2.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R112 m3_4628_86844# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X291 xaa6.xf.XA6.MN0.G xaa6.xf.XA5.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R113 xaa4.xa2.M0.G m3_22620_52900# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X292 xaa3.xa7.MN0.D xaa3.xa6.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R114 li_4836_56708# xaa3.xa1capd.B sky130_fd_pr__res_generic_l1 w=0.44 l=0.36
X293 AVDD PWRUP_1V8 xaa6.xf.XA7.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X294 a_1220_70022# a_788_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R115 AVSS li_6204_61812# sky130_fd_pr__res_generic_l1 w=0.44 l=0.36
X295 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X296 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R116 AVSS m3_37748_96604# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X297 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MP1.G xaa6.xd.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X298 xaa6.xg.XA7.MN2.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X299 xaa5.xa3.xb1_0.G xaa5.xa3.xb2_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R117 m3_4628_100284# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X300 xaa0.xa6.MN0.D xaa0.xa3.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X301 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X302 xaa6.xf.XA5.MN0.G xaa6.xf.XA7.MN1.G xaa6.xf.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X303 a_1220_74698# a_1652_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X304 xaa6.xe.XA1.MN0.D xaa6.xe.XA1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X305 xaa6.xd.XA3.MN0.D xaa6.xd.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X306 xaa6.xg.XA5.MN0.G xaa6.xg.XA3.MN1.G xaa6.xg.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X307 AVDD xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X308 xaa4.xa4.M0.D xaa1.xa3.D xaa4.xa1.M8.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X309 xaa5.xb2_0.MN0.D xaa5.xb1.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X310 xaa0.xa2a.MN0.D xaa0.xa2a.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X311 AVDD PWRUP_1V8 xaa6.xc.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X312 xaa4.xa1.M1.D IBPSR_1U xaa4.xa1.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X313 xaa3.xa8.MP0.D xaa3.xa1b.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X314 xaa5.xa3.xb2_0.D xaa5.xa3.xb1_0.D xaa5.xa3.xc2a.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X315 xaa6.xc.XA5.MN0.G xaa6.xc.XA7.MP1.G xaa6.xc.XA3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X316 xaa6.xd.XA6.MN0.D xaa6.xd.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X317 AVDD xaa4.xa4.M0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X318 xaa5.xa3.xb2_0.G xaa5.xb2_4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X319 xaa1.xa3.D xaa0.xa2a.MN0.D xaa1.xb2.M7.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X320 xaa6.xg.XA7.MP1.G xaa6.xg.XA3.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R118 m3_4628_108924# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R119 AVSS m3_37748_91804# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X321 xaa6.xg.XA4.MN0.D xaa6.xg.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R120 m3_4628_78204# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X322 xaa0.xa1.MN0.G xaa0.xa1.MN2.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X323 xaa3.xa6.MN0.D xaa3.xa5a.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R121 AVSS m3_37748_83164# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X324 xaa6.xc.XA4.MP0.D xaa6.xc.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X325 xaa5.xa4.MN0.D xaa5.xa3.xb1_0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X326 xaa1.xa1.M6.D IBPSR_1U xaa1.xa1.M5.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X327 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MN1.G xaa6.xg.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X328 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MN1.G xaa6.xe.XA7.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X329 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R122 m3_4628_99324# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X330 xaa1.xa3.D PWRUP_1V8 AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X331 xaa6.xg.XA3.MP0.D xaa6.xg.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X332 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X333 xaa0.xa6.MN0.D xaa0.xa3.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X334 xaa1.xa3.D xaa0.xa6.MN0.D xaa1.xa2.M8.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X335 xaa6.xg.XA6.MP0.D xaa6.xg.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X336 xaa6.xe.XA7.MN0.D xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X337 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R123 xaa4.xa2.M0.G m3_22620_61348# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X338 xaa0.xa2a.MN0.D xaa0.xa2a.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X339 xaa1.xa1.M8.D IBPSR_1U xaa1.xa1.M7.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R124 m3_4628_73404# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R125 li_4836_61284# xaa3.xa5a.MN0.D sky130_fd_pr__res_generic_l1 w=0.44 l=0.36
C0 xaa6.xc.XA3.MN0.D a_26092_54158# 0.00176f
C1 xaa6.xf.XA3.MN0.D a_34804_54510# 0.0474f
C2 a_27244_54510# a_28612_54510# 8.89e-19
C3 xaa1.xa4.M0.D m3_37748_103324# 0.111f
C4 li_4468_111644# li_4468_111484# 7.91f
C5 xaa4.xa2.M0.G m3_13044_55188# 0.106f
C6 xaa0.xa2a.MN0.D a_640_59750# 4.85e-19
C7 a_29764_61102# a_29764_60750# 0.0109f
C8 PWRUP_1V8 a_26092_58030# 0.00637f
C9 AVDD a_28612_58030# 0.338f
C10 m2_4468_105884# m3_37668_106204# 0.0138f
C11 a_32284_56974# a_32284_56622# 0.0109f
C12 xaa6.xf.XA7.MP1.G a_34804_56270# 0.1f
C13 xaa6.xf.XA7.MN1.G a_33652_56270# 0.0803f
C14 IBPSR_1U xaa4.xa1.M1.D 0.026f
C15 xaa6.xd.XA1.MN0.G xaa6.xd.XA5.MN0.G 0.00917f
C16 xaa6.xd.XA7.MN0.D xaa6.xd.XA6.MN0.G 3.13e-19
C17 xaa6.xc.XA7.MN1.G a_26092_55918# 7.37e-19
C18 AVDD xaa6.xe.XA3.MN0.D 0.00913f
C19 xaa1.xa4.M0.D m2_4468_78044# 71.5f
C20 xaa6.xe.XA4.MP0.D a_32284_55214# 0.0467f
C21 xaa4.xa2.M0.D xaa4.xa1.M6.D 0.00452f
C22 xaa6.xe.XA5.MN0.G a_31132_54510# 0.00236f
C23 AVDD li_6204_57236# 0.00384f
C24 xaa3.xa5a.MN0.D a_5844_60782# 0.0536f
C25 IBPSR_1U a_640_59750# 0.00137f
C26 xaa5.xa3.xb2_0.G a_26092_60750# 3.06e-19
C27 xaa4.xa2.M0.G a_29764_60750# 1.59e-19
C28 AVDD xaa5.xb2_1.MN0.D 0.543f
C29 PWRUP_1V8 xaa4.xa2.M0.D 0.0181f
C30 xaa0.xa5.MN2.G a_26092_56622# 8.37e-20
C31 xaa6.xe.XA7.MN1.D a_32284_56974# 0.00166f
C32 xaa6.xe.XA1.MN0.G a_31132_56974# 1.06e-19
C33 AVDD a_5844_55502# 0.485f
C34 m2_4468_79004# m3_37748_79324# 0.0138f
C35 xaa6.xg.XA5.MN0.D xaa6.xg.XA5.MN0.G 0.109f
C36 xaa6.xd.XA1.MN0.G a_28612_53102# 0.0658f
C37 xaa6.xd.XA7.MN1.D a_29764_53102# 8.73e-21
C38 a_37324_55918# a_37324_55566# 0.0109f
C39 xaa1.xa4.M0.D m1_4468_92444# 67.7f
C40 xaa6.xg.XA7.MN1.D a_37324_53454# 6.39e-19
C41 xaa6.xf.XA7.MP1.G a_34804_53806# 0.00375f
C42 xaa6.xf.XA7.MN1.G a_33652_53806# 0.113f
C43 xaa1.xa4.M0.D m3_4788_86844# 0.0138f
C44 a_27244_53806# a_28612_53806# 8.89e-19
C45 li_4468_95164# li_4468_94364# 39.3f
C46 xaa1.xa2.M6.D xaa1.xa2.M5.D 0.0488f
C47 xaa4.xa2.M0.G a_28612_63214# 0.0361f
C48 xaa5.xb1.MN1.G xaa5.xb2_3.MN0.D 0.04f
C49 xbb0.xa1.XA1.N a_788_72222# 7.07e-19
C50 a_26092_58030# a_26092_57678# 0.0109f
C51 xaa0.xa2a.MN0.D a_244_56622# 2.1e-19
C52 a_32284_58030# xaa6.xe.XA7.MN1.D 0.0658f
C53 a_31132_58030# xaa6.xe.XA1.MN0.G 1.35e-19
C54 PWRUP_1V8 xaa6.xg.XA7.MN2.D 0.0119f
C55 AVDD a_27244_56974# 0.405f
C56 m2_4468_92444# m3_37668_92764# 0.0138f
C57 PWRUP_1V8 a_34804_53454# 0.0705f
C58 xaa6.xc.XA7.MN1.G a_28612_54862# 7.1e-20
C59 xaa6.xc.XA7.MP1.G a_27244_54862# 0.097f
C60 a_29764_56622# xaa6.xd.XA5.MN0.G 6.14e-19
C61 xaa6.xf.XA6.MP0.D a_33652_56270# 0.0467f
C62 xaa6.xc.XA7.MN1.D a_26092_54510# 0.0736f
C63 xaa6.xe.XA1.MN0.G xaa6.xf.XA3.MP0.D 0.00218f
C64 AVDD a_37324_53454# 0.369f
C65 xaa6.xf.XA3.MP0.D a_34804_54510# 2.16e-19
C66 xaa6.xf.XA3.MN0.D a_33652_54510# 2.16e-19
C67 xaa1.xa4.M0.D m3_37668_103324# 0.074f
C68 xaa4.xa2.M0.G m3_22620_56068# 0.0273f
C69 li_4468_78044# m1_4468_78044# 23f
C70 xaa0.xa2a.MN0.D a_n908_59750# 7.26e-19
C71 a_4692_60430# a_5844_60430# 0.00133f
C72 AVDD a_27244_58030# 0.343f
C73 xaa0.xa5.MN0.D xaa0.xa1.MN2.S 0.00385f
C74 xaa6.xf.XA7.MP1.G a_33652_56270# 0.0268f
C75 xaa6.xf.XA7.MN1.G a_32284_56270# 7.1e-20
C76 xaa6.xd.XA7.MN1.D xaa6.xd.XA5.MN0.G 0.29f
C77 xaa6.xd.XA7.MN1.G xaa6.xd.XA6.MN0.G 0.329f
C78 AVDD xaa6.xd.XA3.MN0.D 0.00913f
C79 xaa1.xa4.M0.D m2_4468_79004# 71.5f
C80 xaa4.xa2.M0.D a_11712_54334# 0.151f
C81 AVDD li_6132_57236# 0.00142f
C82 a_32284_53102# a_33652_53102# 8.89e-19
C83 li_4468_78044# li_4468_77884# 7.91f
C84 xaa3.xa5a.MN0.D a_4692_60782# 0.0583f
C85 a_29764_62510# PWRUP_1V8 1.55e-20
C86 IBPSR_1U a_n908_59750# 0.0719f
C87 xaa4.xa2.M0.G a_28612_60750# 0.0273f
C88 a_28612_62158# a_28612_61806# 0.0109f
C89 AVDD xaa5.xa3.xb1_0.D 1.88f
C90 xaa6.xe.XA7.MN0.D a_32284_57326# 0.0525f
C91 xaa6.xe.XA7.MN1.D a_31132_56974# 0.0092f
C92 xaa6.xd.XA1.MN0.G a_32284_56974# 0.0725f
C93 AVDD a_4692_55502# 0.00171f
C94 m2_4468_79004# m3_37668_79324# 0.0138f
C95 xaa6.xf.XA1.MN0.G a_37324_53454# 1.11e-19
C96 xaa6.xc.XA5.MN0.G a_27244_55566# 0.0889f
C97 xaa6.xc.XA6.MN0.G xaa6.xc.XA4.MP0.D 0.0357f
C98 xaa6.xf.XA5.MN0.G xaa6.xg.XA5.MN0.G 0.00217f
C99 xaa6.xd.XA7.MN1.D a_28612_53102# 5.24e-20
C100 xaa1.xa4.M0.D m1_4468_93404# 67.7f
C101 xaa6.xf.XA7.MP1.G a_33652_53806# 0.00282f
C102 xaa6.xf.XA7.MN1.G a_32284_53806# 7.1e-20
C103 xaa1.xa4.M0.D m3_4628_86844# 0.0276f
C104 xaa6.xg.XA3.MN1.G a_37324_53102# 0.00349f
C105 a_4692_63070# a_4692_62718# 0.0109f
C106 xaa5.xb1.MN1.G a_29764_63214# 0.00504f
C107 xaa4.xa2.M0.G a_27244_63214# 6.72e-19
C108 a_788_76898# a_2948_74698# 2.35e-20
C109 m1_4468_105884# m2_4468_105884# 12.9f
C110 a_31132_58030# xaa6.xe.XA7.MN1.D 0.0711f
C111 PWRUP_1V8 xaa6.xg.XA7.MN0.G 0.077f
C112 xaa1.xa3.D xaa4.xa1.M8.D 0.0639f
C113 a_32284_58030# xaa6.xd.XA1.MN0.G 0.0342f
C114 AVDD a_26092_56974# 0.00159f
C115 xaa1.xa4.M0.D li_4468_85564# 23f
C116 a_36172_56974# xaa6.xg.XA5.MN0.G 1.67e-19
C117 xaa6.xe.XA7.MP1.G a_32284_55214# 0.027f
C118 xaa6.xe.XA7.MN1.G a_33652_55214# 7.1e-20
C119 PWRUP_1V8 a_33652_53454# 0.0658f
C120 xaa6.xc.XA7.MN1.G a_27244_54862# 0.00608f
C121 xaa6.xc.XA7.MP1.G a_26092_54862# 0.029f
C122 a_26092_56270# a_27244_56270# 0.00133f
C123 xaa6.xc.XA6.MP0.D xaa6.xc.XA6.MN0.G 0.0116f
C124 CK a_37324_52750# 0.00287f
C125 xaa6.xe.XA1.MN0.G xaa6.xe.XA3.MP0.D 0.00238f
C126 AVDD a_36172_53454# 0.00151f
C127 xaa6.xf.XA3.MP0.D a_33652_54510# 0.0467f
C128 a_26092_54510# a_27244_54510# 0.00133f
C129 a_10092_54510# xaa4.xa1.M5.D 2.99e-19
C130 xaa1.xa4.M0.D m3_4788_104124# 0.0138f
C131 li_4468_112444# li_4468_111644# 39.3f
C132 xaa4.xa2.M0.G m3_22548_56068# 0.0137f
C133 xaa1.xa1.M5.D a_n908_59750# 8.62e-20
C134 xaa1.xb2.M0.D a_640_60278# 0.00155f
C135 xaa3.xa4.MN0.D a_5844_60430# 0.0897f
C136 a_28612_61102# a_28612_60750# 0.0109f
C137 xaa1.xa1.M2.D xaa1.xa1.M1.D 0.0488f
C138 AVDD a_26092_58030# 0.00527f
C139 a_31132_56974# a_31132_56622# 0.0109f
C140 xaa6.xc.XA1.MN0.G xaa6.xd.XA5.MN0.G 0.00881f
C141 xaa6.xd.XA7.MP1.G xaa6.xd.XA6.MN0.G 0.524f
C142 xaa6.xd.XA7.MN1.G xaa6.xc.XA6.MN0.G 3.47e-19
C143 a_11712_57502# a_11712_55918# 0.00223f
C144 AVDD xaa6.xd.XA3.MP0.D 0.133f
C145 xaa1.xa4.M0.D m2_4468_79964# 71.5f
C146 xaa6.xg.XA5.MN0.G xaa6.xg.XA3.MP0.D 0.0488f
C147 xaa6.xe.XA4.MN0.D a_31132_55214# 0.0472f
C148 xaa4.xa2.M0.D xaa4.xa1.M7.D 0.00653f
C149 xaa6.xd.XA5.MN0.G a_29764_54510# 0.00236f
C150 li_4468_101084# m1_4468_101084# 23f
C151 xaa5.xa3.xb1_0.D xaa5.xb1.MN1.D 0.00329f
C152 IBPSR_1U xaa4.xa4.M0.D 0.00246f
C153 xaa5.xb1.MN1.G a_29764_60750# 0.00139f
C154 xaa4.xa2.M0.G a_27244_60750# 3.15e-19
C155 xaa1.xa2.M2.D a_n908_61510# 2.99e-19
C156 xaa1.xa2.M1.D xaa1.xa2.M0.D 0.0488f
C157 AVDD xaa5.xa4.MN0.D 0.227f
C158 m1_4468_72284# m2_4468_72284# 12.9f
C159 PWRUP_1V8 a_36172_55918# 0.00682f
C160 xaa6.xe.XA7.MN0.D a_31132_57326# 0.055f
C161 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MN2.D 0.0372f
C162 xaa6.xe.XA7.MN1.D a_29764_56974# 1.31e-19
C163 xaa6.xg.XA7.MP1.G xaa6.xg.XA7.MN0.D 0.117f
C164 xaa6.xd.XA1.MN0.G a_31132_56974# 0.0672f
C165 xaa6.xe.XA7.MP1.G a_32284_57326# 0.0964f
C166 AVDD xaa4.xa2.M0.D 7.31f
C167 xaa6.xf.XA1.MN0.G a_36172_53454# 0.00212f
C168 xaa6.xc.XA5.MN0.G a_26092_55566# 0.112f
C169 xaa6.xc.XA6.MN0.G xaa6.xc.XA4.MN0.D 0.0093f
C170 a_36172_55918# a_36172_55566# 0.0109f
C171 xaa1.xa4.M0.D m1_4468_94364# 67.7f
C172 xaa1.xa4.M0.D m3_37748_87004# 0.111f
C173 xaa6.xg.XA3.MN1.G a_36172_53102# 7.28e-19
C174 a_26092_53806# a_27244_53806# 0.00133f
C175 li_4468_95324# li_4468_95164# 7.91f
C176 a_5844_63070# xaa3.xa6.MN0.D 0.0658f
C177 xaa5.xa3.xb1_0.G a_27244_63214# 0.00131f
C178 xaa5.xb1.MN1.G a_28612_63214# 9.6e-19
C179 xaa0.xa2a.MN0.D xaa0.xa3.MN1.G 0.00708f
C180 PWRUP_1V8 xaa6.xf.XA7.MN2.D 0.0119f
C181 a_31132_58030# xaa6.xd.XA1.MN0.G 0.0408f
C182 xaa4.xa4.M0.D a_11712_57502# 0.154f
C183 AVDD xaa6.xg.XA7.MN2.D 0.00837f
C184 PWRUP_1V8 a_32284_53454# 0.0674f
C185 xaa6.xe.XA7.MP1.G a_31132_55214# 0.0944f
C186 xaa6.xe.XA7.MN1.G a_32284_55214# 0.0761f
C187 xaa6.xc.XA7.MN1.G a_26092_54862# 0.0724f
C188 xaa6.xe.XA6.MP0.D a_32284_56270# 0.0467f
C189 xaa6.xc.XA6.MN0.D xaa6.xc.XA6.MN0.G 0.0093f
C190 CK a_36172_52750# 0.00871f
C191 xaa6.xe.XA7.MN1.D xaa6.xe.XA3.MP0.D 0.0844f
C192 xaa6.xe.XA1.MN0.G xaa6.xe.XA3.MN0.D 6.01e-19
C193 xaa6.xg.XA7.MP1.G xaa6.xg.XA4.MP0.D 0.0615f
C194 AVDD a_34804_53454# 0.00151f
C195 a_10092_54510# xaa4.xa1.M6.D 5.84e-19
C196 xaa1.xa4.M0.D m3_4628_104124# 0.0276f
C197 xaa4.xa2.M0.G m3_13116_56244# 0.0634f
C198 xaa3.xa4.MN0.D a_4692_60430# 0.117f
C199 PWRUP_1V8 xaa3.xa1capd.B 0.00221f
C200 AVDD a_5844_57790# 0.364f
C201 xaa0.xa5.MN0.D a_n908_55214# 3.18e-19
C202 xaa6.xg.XA7.MN2.D a_36172_56622# 0.00176f
C203 a_36172_56974# a_37324_56974# 0.00133f
C204 xaa6.xc.XA1.MN0.G xaa6.xc.XA5.MN0.G 0.01f
C205 xaa6.xg.XA7.MN1.D a_37324_55918# 0.00149f
C206 AVDD xaa6.xc.XA3.MP0.D 0.133f
C207 xaa1.xa4.M0.D m2_4468_80924# 71.5f
C208 xaa6.xg.XA5.MN0.G xaa6.xg.XA3.MN0.D 0.0488f
C209 xaa6.xd.XA5.MN0.G a_28612_54510# 0.00224f
C210 xaa4.xa1.M0.D a_10092_52750# 0.00155f
C211 a_31132_53102# a_32284_53102# 0.00133f
C212 xbb1.xa3.M4.D xbb1.xa3.M3.D 0.0488f
C213 li_4468_78844# li_4468_78044# 39.3f
C214 a_27244_62158# a_27244_61806# 0.0109f
C215 CK a_29764_61454# 3.97e-20
C216 AVDD a_29764_62510# 0.00139f
C217 PWRUP_1V8 a_34804_55918# 0.00684f
C218 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MN0.G 0.0363f
C219 xaa6.xg.XA7.MN1.G xaa6.xg.XA7.MN0.D 0.0449f
C220 xaa6.xd.XA1.MN0.G a_29764_56974# 0.00134f
C221 xaa6.xd.XA7.MN1.D a_31132_56974# 1.31e-19
C222 xaa6.xe.XA7.MP1.G a_31132_57326# 9.02e-20
C223 xaa6.xe.XA7.MN1.G a_32284_57326# 0.00174f
C224 AVDD a_37324_55918# 0.386f
C225 xaa6.xf.XA1.MN0.G a_34804_53454# 0.0733f
C226 xaa6.xc.XA1.MN0.G a_27244_53102# 0.0711f
C227 xaa1.xa4.M0.D m1_4468_95324# 67.7f
C228 xaa1.xa4.M0.D m3_37668_87004# 0.074f
C229 a_37324_57678# m1_37504_57930# 0.0182f
C230 a_4692_63070# xaa3.xa6.MN0.D 0.0732f
C231 xaa5.xa3.xb1_0.G a_26092_63214# 0.00428f
C232 a_788_76898# xaa1.xa4.M0.D 0.0454f
C233 m1_4468_106844# m2_4468_106844# 12.9f
C234 xaa0.xa2a.MN0.D a_244_56974# 3.94e-19
C235 a_36172_58030# a_37324_58030# 0.00133f
C236 PWRUP_1V8 xaa6.xe.XA7.MN2.D 0.0119f
C237 a_29764_58030# xaa6.xd.XA1.MN0.G 0.00237f
C238 AVDD xaa6.xg.XA7.MN0.G 0.479f
C239 PWRUP_1V8 a_31132_53454# 0.0689f
C240 xaa1.xa4.M0.D li_4468_86524# 23f
C241 xaa6.xe.XA7.MN1.G a_31132_55214# 0.00134f
C242 xaa6.xe.XA6.MN0.D a_32284_56270# 2.16e-19
C243 xaa6.xe.XA6.MP0.D a_31132_56270# 2.16e-19
C244 CK a_34804_52750# 0.00126f
C245 xaa6.xe.XA7.MN1.D xaa6.xe.XA3.MN0.D 0.0425f
C246 xaa6.xg.XA7.MP1.G xaa6.xg.XA4.MN0.D 0.056f
C247 xaa6.xg.XA7.MN1.G xaa6.xg.XA4.MP0.D 1.09e-19
C248 xaa6.xd.XA1.MN0.G xaa6.xe.XA3.MP0.D 2.36e-19
C249 AVDD a_33652_53454# 0.368f
C250 xaa6.xe.XA3.MP0.D a_32284_54510# 0.0467f
C251 xaa1.xa4.M0.D m3_37748_104284# 0.111f
C252 li_4468_112604# li_4468_112444# 7.91f
C253 xaa4.xa2.M0.G m3_13044_56244# 0.106f
C254 xaa1.xa3.D a_2948_70022# 0.201f
C255 li_4468_79004# m1_4468_79004# 23f
C256 a_27244_61102# a_27244_60750# 0.0109f
C257 xaa0.xa6.MN0.D a_244_56270# 0.00172f
C258 AVDD a_4692_57790# 0.00171f
C259 m2_4468_106844# m3_37748_107164# 0.0138f
C260 xaa0.xa3.MN1.G xaa0.xa1.MN2.S 0.0608f
C261 xaa6.xf.XA1.MN0.G a_37324_55918# 1.11e-19
C262 xaa6.xe.XA7.MP1.G a_32284_56270# 0.0268f
C263 xaa6.xe.XA7.MN1.G a_33652_56270# 7.1e-20
C264 a_29764_56974# a_29764_56622# 0.0109f
C265 xaa6.xc.XA7.MN1.D xaa6.xc.XA5.MN0.G 0.29f
C266 xaa6.xc.XA7.MN0.D xaa6.xc.XA6.MN0.G 3.13e-19
C267 xaa6.xg.XA7.MN1.D a_36172_55918# 0.00829f
C268 xaa6.xg.XA7.MP1.G xaa6.xg.XA6.MP0.D 0.0619f
C269 AVDD xaa6.xc.XA3.MN0.D 0.00913f
C270 xaa1.xa4.M0.D m2_4468_81884# 71.5f
C271 xaa6.xg.XA4.MP1.G xaa6.xg.XA4.MP0.D 0.0093f
C272 xaa6.xd.XA4.MN0.D a_29764_55214# 0.0472f
C273 xaa6.xg.XA5.MN0.G xaa6.xg.XA3.MN1.G 0.0308f
C274 AVDD li_6204_59524# 0.00384f
C275 xaa5.xa3.xb2_0.D a_27244_61454# 0.0972f
C276 xaa5.xb2_1.MN0.D a_29764_61806# 0.00263f
C277 xaa5.xa3.xb1_0.G a_26092_60750# 0.0733f
C278 a_29764_62158# xaa5.xb2_0.MN0.D 0.0682f
C279 AVDD a_28612_62510# 0.352f
C280 m1_4468_73244# m2_4468_73244# 12.9f
C281 xaa6.xg.XA7.MN1.G xaa6.xg.XA7.MP1.G 0.141f
C282 xaa6.xf.XA1.MN0.G xaa6.xg.XA7.MN0.G 0.00299f
C283 xaa6.xd.XA7.MN1.D a_29764_56974# 0.0092f
C284 xaa6.xe.XA7.MN1.G a_31132_57326# 0.0781f
C285 AVDD a_36172_55918# 0.00151f
C286 xaa6.xf.XA1.MN0.G a_33652_53454# 0.0676f
C287 xaa6.xc.XA7.MN1.D a_27244_53102# 5.24e-20
C288 a_10092_55566# xaa4.xa1.M8.D 0.0223f
C289 xaa6.xc.XA1.MN0.G a_26092_53102# 0.0727f
C290 xaa6.xe.XA7.MN1.G a_33652_53806# 7.1e-20
C291 xaa6.xe.XA7.MP1.G a_32284_53806# 0.00282f
C292 xaa6.xe.XA5.MN0.G xaa6.xf.XA5.MN0.G 0.00217f
C293 a_34804_55918# a_34804_55566# 0.0109f
C294 xaa1.xa4.M0.D m1_4468_96284# 67.7f
C295 xaa6.xc.XA7.MN1.G xaa6.xc.XA1.MN0.D 0.123f
C296 a_36172_57678# m1_37504_57930# 6.53e-19
C297 xaa1.xa4.M0.D m3_4788_87804# 0.0138f
C298 li_4468_96124# li_4468_95324# 39.3f
C299 xbb0.xa1.XA1.N a_n76_72222# 0.113f
C300 xaa0.xa2a.MN0.D a_n908_56974# 3.79e-19
C301 PWRUP_1V8 xaa6.xd.XA7.MN2.D 0.0119f
C302 a_29764_58030# xaa6.xd.XA7.MN1.D 0.0693f
C303 AVDD xaa6.xf.XA7.MN2.D 0.00837f
C304 m2_4468_93404# m3_37748_93724# 0.0138f
C305 PWRUP_1V8 a_29764_53454# 0.0705f
C306 xaa0.xa5.MN0.D a_n908_54510# 3.3e-20
C307 a_26092_56622# xaa6.xc.XA5.MN0.G 6.14e-19
C308 xaa6.xe.XA6.MN0.D a_31132_56270# 0.0474f
C309 xaa6.xg.XA7.MP1.G xaa6.xg.XA4.MP1.G 0.0436f
C310 a_34804_56974# xaa6.xf.XA5.MN0.G 1.55e-19
C311 xaa6.xg.XA7.MN1.G xaa6.xg.XA4.MN0.D 1.09e-19
C312 xaa6.xd.XA1.MN0.G xaa6.xe.XA3.MN0.D 0.00287f
C313 AVDD a_32284_53454# 0.367f
C314 xaa4.xa2.M0.D a_11712_52750# 0.0717f
C315 a_10092_54510# xaa4.xa1.M7.D 0.00155f
C316 xaa6.xe.XA3.MN0.D a_32284_54510# 2.16e-19
C317 xaa6.xe.XA3.MP0.D a_31132_54510# 2.16e-19
C318 xaa1.xa4.M0.D m3_37668_104284# 0.074f
C319 xaa4.xa2.M0.G m3_22620_57124# 0.0273f
C320 a_2084_70022# a_2948_70022# 0.00813f
C321 a_5844_60782# a_5844_60430# 0.0109f
C322 xaa0.xa6.MN0.D a_n908_56270# 3.59e-19
C323 AVDD xaa3.xa1capd.B 1.12f
C324 m2_4468_106844# m3_37668_107164# 0.0138f
C325 a_n908_56270# xaa0.xa1.MN0.G 1.72e-19
C326 a_244_56270# a_244_55918# 0.0109f
C327 a_34804_56974# a_36172_56974# 8.89e-19
C328 xaa0.xa5.MN0.D a_244_55566# 1.28e-19
C329 xaa0.xa3.MN1.G a_244_55214# 0.0674f
C330 xaa6.xe.XA7.MP1.G a_31132_56270# 0.0985f
C331 xaa6.xe.XA7.MN1.G a_32284_56270# 0.0819f
C332 xaa6.xf.XA1.MN0.G a_36172_55918# 0.00205f
C333 xaa6.xc.XA7.MN1.G xaa6.xd.XA6.MN0.G 3.47e-19
C334 xaa6.xc.XA7.MP1.G xaa6.xc.XA6.MN0.G 0.524f
C335 xaa0.xa5.MN2.G xaa6.xc.XA5.MN0.G 9.76e-20
C336 xaa3.xa1b.MN0.D xbb1.xa3.M6.D 1.38e-19
C337 PWRUP_1V8 a_36172_54862# 0.00561f
C338 xaa6.xg.XA7.MP1.G xaa6.xg.XA6.MN0.D 0.056f
C339 xaa6.xg.XA7.MN1.G xaa6.xg.XA6.MP0.D 0.0287f
C340 AVDD a_10092_54510# 0.0011f
C341 xaa1.xa4.M0.D m2_4468_82844# 71.5f
C342 xaa6.xc.XA5.MN0.G a_27244_54510# 0.00224f
C343 AVDD li_6132_59524# 0.00142f
C344 a_29764_53102# a_31132_53102# 8.89e-19
C345 li_4468_102044# m1_4468_102044# 23f
C346 li_4468_79004# li_4468_78844# 7.91f
C347 xaa5.xa3.xb2_0.D a_26092_61454# 0.00277f
C348 xaa5.xb2_1.MN0.D a_28612_61806# 0.00224f
C349 a_26092_62158# a_26092_61806# 0.0109f
C350 a_28612_62158# xaa5.xb2_0.MN0.D 0.0674f
C351 AVDD a_27244_62510# 0.388f
C352 xaa6.xf.XA7.MN1.D xaa6.xg.XA7.MN0.G 2.06e-19
C353 xaa6.xd.XA7.MN1.D a_28612_56974# 0.00166f
C354 xaa6.xc.XA1.MN0.G a_29764_56974# 0.0677f
C355 AVDD a_34804_55918# 0.00151f
C356 m2_4468_79964# m3_37748_80284# 0.0138f
C357 xaa6.xe.XA1.MN0.G a_34804_53454# 1.02e-19
C358 xaa6.xf.XA7.MN1.D a_33652_53454# 6.39e-19
C359 xaa6.xc.XA7.MN1.D a_26092_53102# 8.73e-21
C360 xaa6.xe.XA7.MP1.G a_31132_53806# 0.00375f
C361 xaa6.xe.XA7.MN1.G a_32284_53806# 0.115f
C362 xaa1.xa4.M0.D m1_4468_97244# 67.7f
C363 xaa1.xa4.M0.D m3_4628_87804# 0.0276f
C364 xaa1.xa3.D xaa1.xa2.M1.D 7.7e-19
C365 xaa1.xa2.M7.D xaa1.xa2.M6.D 0.0488f
C366 a_4692_63070# a_5844_63070# 0.00133f
C367 m1_4468_107804# m2_4468_107804# 12.9f
C368 a_34804_58030# a_36172_58030# 8.89e-19
C369 PWRUP_1V8 xaa6.xc.XA7.MN2.D 0.0123f
C370 a_29764_58030# xaa6.xc.XA1.MN0.G 0.0354f
C371 a_28612_58030# xaa6.xd.XA7.MN1.D 0.0674f
C372 AVDD xaa6.xe.XA7.MN2.D 0.00837f
C373 m2_4468_93404# m3_37668_93724# 0.0138f
C374 xaa6.xg.XA7.MN1.D a_37324_54862# 0.00464f
C375 PWRUP_1V8 a_28612_53454# 0.0658f
C376 xaa1.xa4.M0.D li_4468_87484# 23f
C377 xaa6.xg.XA6.MN0.D xaa6.xg.XA6.MP0.D 0.00918f
C378 xaa6.xg.XA7.MN1.G xaa6.xg.XA4.MP1.G 0.0438f
C379 xaa6.xd.XA1.MN0.G xaa6.xd.XA3.MN0.D 0.00303f
C380 xaa0.xa5.MN0.D xaa0.xa2a.MN0.G 7.05e-20
C381 AVDD a_31132_53454# 0.00151f
C382 xaa6.xe.XA3.MN0.D a_31132_54510# 0.0474f
C383 xaa6.xg.XA3.MN0.D xaa6.xg.XA3.MP0.D 0.00918f
C384 xaa1.xa4.M0.D m3_4788_105084# 0.0138f
C385 li_4468_113404# li_4468_112604# 39.3f
C386 xaa4.xa2.M0.G m3_22548_57124# 0.0137f
C387 a_26092_61102# a_26092_60750# 0.0109f
C388 xaa5.xb1.MN0.D a_29764_60750# 0.00176f
C389 xaa1.xa1.M6.D a_n908_59750# 6.46e-20
C390 a_640_60806# a_640_60278# 0.00702f
C391 xaa0.xa6.MN0.D xaa0.xa5.MN2.D 3.31e-19
C392 AVDD a_5844_58142# 0.388f
C393 xaa0.xa5.MN2.D xaa0.xa1.MN0.G 2.29e-19
C394 a_28612_56974# a_28612_56622# 0.0109f
C395 xaa6.xf.XA7.MN2.D a_34804_56622# 0.00176f
C396 xaa0.xa3.MN1.G a_n908_55214# 0.0661f
C397 xaa6.xe.XA7.MN1.G a_31132_56270# 0.00344f
C398 xaa6.xf.XA1.MN0.G a_34804_55918# 0.00217f
C399 xaa6.xc.XA7.MN1.G xaa6.xc.XA6.MN0.G 0.329f
C400 IBPSR_1U xbb1.xa3.M6.D 0.0484f
C401 PWRUP_1V8 a_34804_54862# 0.00561f
C402 xaa0.xa5.MN0.D a_n908_55566# 0.00385f
C403 xaa6.xg.XA7.MN1.G xaa6.xg.XA6.MN0.D 0.0158f
C404 AVDD a_37324_54862# 0.382f
C405 xaa1.xa4.M0.D m2_4468_83804# 71.5f
C406 xaa6.xd.XA4.MP0.D a_28612_55214# 0.0467f
C407 xaa6.xc.XA5.MN0.G a_26092_54510# 0.00236f
C408 xbb1.xa3.M6.D a_4308_51918# 6.46e-20
C409 a_37324_53454# a_37324_53102# 0.0109f
C410 CK a_26092_61454# 7.25e-20
C411 xaa5.xa3.xb2_0.D PWRUP_1V8 0.00217f
C412 xaa5.xa3.xb1_0.D a_28612_61806# 4.81e-19
C413 AVDD a_26092_62510# 0.00173f
C414 m1_4468_74204# m2_4468_74204# 12.9f
C415 PWRUP_1V8 a_31132_55918# 0.00682f
C416 xaa6.xe.XA1.MN0.G xaa6.xg.XA7.MN0.G 0.00217f
C417 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MN2.D 0.0372f
C418 xaa6.xd.XA7.MN0.D a_29764_57326# 0.055f
C419 xaa6.xc.XA1.MN0.G a_28612_56974# 0.0736f
C420 AVDD a_33652_55918# 0.385f
C421 m2_4468_79964# m3_37668_80284# 0.0138f
C422 xaa6.xd.XA5.MN0.G xaa6.xe.XA5.MN0.G 0.00217f
C423 xaa6.xe.XA1.MN0.G a_33652_53454# 0.00209f
C424 xaa6.xe.XA7.MN1.G a_31132_53806# 0.114f
C425 a_33652_55918# a_33652_55566# 0.0109f
C426 xaa1.xa4.M0.D m1_4468_98204# 67.7f
C427 xaa1.xa4.M0.D m3_37748_87964# 0.111f
C428 a_37324_54158# a_37324_53806# 0.0109f
C429 li_4468_96284# li_4468_96124# 7.91f
C430 a_28612_58030# xaa6.xc.XA1.MN0.G 0.0493f
C431 AVDD xaa6.xd.XA7.MN2.D 0.00837f
C432 xaa6.xg.XA7.MN1.D a_36172_54862# 0.00652f
C433 PWRUP_1V8 a_27244_53454# 0.0674f
C434 xaa6.xd.XA6.MN0.D a_29764_56270# 0.0474f
C435 xaa6.xf.XA1.MN0.G a_37324_54862# 1.11e-19
C436 xaa6.xd.XA7.MN1.G a_29764_55214# 0.00134f
C437 xaa6.xd.XA7.MN1.D xaa6.xd.XA3.MN0.D 0.0425f
C438 xaa6.xd.XA1.MN0.G xaa6.xd.XA3.MP0.D 3.58e-19
C439 AVDD a_29764_53454# 0.00151f
C440 a_37324_54862# a_37324_54510# 0.0109f
C441 xaa6.xg.XA3.MN1.G xaa6.xg.XA3.MP0.D 9.89e-20
C442 xaa1.xa4.M0.D m3_4628_105084# 0.0276f
C443 xaa4.xa2.M0.G m3_13116_57300# 0.0634f
C444 a_2084_70022# xaa1.xa3.D 0.0226f
C445 li_4468_79964# m1_4468_79964# 23f
C446 a_5844_60782# xaa3.xa4.MN0.D 0.0658f
C447 a_4692_60782# a_4692_60430# 0.0109f
C448 xaa0.xa6.MN0.D xaa0.xa5.MN0.D 0.01f
C449 AVDD a_4692_58142# 0.00171f
C450 a_n908_56270# a_n908_55918# 0.0109f
C451 a_244_56270# xaa0.xa5.MP1.D 0.00176f
C452 a_33652_56974# a_34804_56974# 0.00133f
C453 xaa0.xa5.MN0.D xaa0.xa1.MN0.G 0.15f
C454 xaa0.xa3.MN1.G xaa0.xa3.MP0.D 0.00991f
C455 xaa6.xf.XA1.MN0.G a_33652_55918# 1.35e-19
C456 xaa6.xf.XA7.MN1.D a_34804_55918# 0.00829f
C457 IBPSR_1U xaa4.xa1.M2.D 0.026f
C458 AVDD a_36172_54862# 0.00151f
C459 xaa1.xa4.M0.D m2_4468_84764# 71.5f
C460 xaa6.xf.XA5.MN0.G xaa6.xf.XA3.MN0.D 0.0488f
C461 a_28612_53102# a_29764_53102# 0.00133f
C462 li_4468_79804# li_4468_79004# 39.3f
C463 AVDD xaa5.xb2_2.MN0.D 0.543f
C464 CK PWRUP_1V8 0.31f
C465 xaa5.xa3.xb1_0.D a_27244_61806# 0.154f
C466 a_27244_62158# xaa5.xa3.xc2a.D 0.00176f
C467 PWRUP_1V8 a_29764_55918# 0.00684f
C468 a_37324_57678# a_37324_57326# 0.0109f
C469 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN2.D 0.0101f
C470 xaa6.xd.XA7.MN0.D a_28612_57326# 0.0525f
C471 xaa6.xd.XA7.MN1.G a_29764_57326# 0.0797f
C472 xaa6.xc.XA1.MN0.G a_27244_56974# 0.00218f
C473 xaa6.xf.XA7.MP1.G xaa6.xg.XA7.MP1.G 0.00435f
C474 xaa6.xf.XA7.MN1.G xaa6.xg.XA7.MN1.G 0.00646f
C475 AVDD a_32284_55918# 0.385f
C476 xaa6.xe.XA1.MN0.G a_32284_53454# 0.0739f
C477 xaa1.xa4.M0.D m1_4468_99164# 67.7f
C478 xaa1.xa4.M0.D m3_37668_87964# 0.074f
C479 xaa3.xa1b.MN0.D a_4692_62366# 0.0046f
C480 a_788_76898# a_1652_76898# 0.107f
C481 xbb0.xa1.XA1.N a_n940_70022# 0.0295f
C482 a_n76_76898# xaa1.xa4.M0.D 0.0448f
C483 m1_4468_108764# m2_4468_108764# 12.9f
C484 a_33652_58030# a_34804_58030# 0.00133f
C485 PWRUP_1V8 a_n908_56270# 6.76e-19
C486 a_27244_58030# xaa6.xc.XA1.MN0.G 0.0026f
C487 AVDD xaa6.xc.XA7.MN2.D 0.00837f
C488 PWRUP_1V8 a_26092_53454# 0.0693f
C489 xaa1.xa4.M0.D li_4468_88444# 23f
C490 xaa6.xd.XA6.MP0.D a_29764_56270# 2.16e-19
C491 xaa6.xd.XA6.MN0.D a_28612_56270# 2.16e-19
C492 xaa6.xf.XA1.MN0.G a_36172_54862# 0.00205f
C493 xaa6.xd.XA7.MP1.G a_29764_55214# 0.096f
C494 xaa6.xd.XA7.MN1.G a_28612_55214# 0.0745f
C495 xaa6.xd.XA7.MN1.D xaa6.xd.XA3.MP0.D 0.0844f
C496 xaa6.xc.XA1.MN0.G xaa6.xd.XA3.MN0.D 3.2e-19
C497 xaa0.xa5.MN0.D a_n908_54862# 6.02e-20
C498 AVDD a_28612_53454# 0.368f
C499 xaa6.xd.XA3.MN0.D a_29764_54510# 0.0474f
C500 xaa6.xg.XA3.MN1.G xaa6.xg.XA3.MN0.D 0.0288f
C501 xaa1.xa4.M0.D m3_37748_105244# 0.111f
C502 li_4468_113564# li_4468_113404# 7.91f
C503 xaa4.xa2.M0.G m3_13044_57300# 0.106f
C504 a_1652_72222# a_2948_70022# 0.00121f
C505 a_4692_60782# xaa3.xa4.MN0.D 0.0728f
C506 xaa1.xb2.M7.D a_640_60278# 5.84e-19
C507 xaa0.xa6.MN0.D a_244_56622# 0.00581f
C508 AVDD xaa3.xa2.MN0.D 0.72f
C509 a_27244_56974# a_27244_56622# 0.0109f
C510 xaa0.xa5.MN2.D a_n908_55918# 0.00176f
C511 xaa0.xa5.MN0.D a_244_55918# 0.00328f
C512 xaa0.xa3.MN1.G a_244_55566# 0.0665f
C513 xaa6.xe.XA1.MN0.G a_34804_55918# 1.02e-19
C514 xaa6.xf.XA7.MN1.D a_33652_55918# 0.00149f
C515 AVDD a_34804_54862# 0.00151f
C516 xaa1.xa4.M0.D m2_4468_85724# 71.5f
C517 xaa6.xc.XA4.MP0.D a_27244_55214# 0.0467f
C518 xaa6.xf.XA5.MN0.G xaa6.xf.XA3.MP0.D 0.0488f
C519 AVDD li_6204_61812# 0.00384f
C520 a_36172_53454# a_36172_53102# 0.0109f
C521 li_4468_103004# m1_4468_103004# 23f
C522 xaa0.xa6.MN0.D a_n908_59750# 7.06e-19
C523 xaa5.xa3.xb1_0.D a_26092_61806# 0.0147f
C524 xaa3.xa1b.MN0.D a_4692_60078# 0.00455f
C525 a_28612_62158# a_29764_62158# 0.00133f
C526 AVDD xaa5.xa3.xb2_0.D 1.82f
C527 m1_4468_75164# m2_4468_75164# 12.9f
C528 xaa6.xc.XA7.MN1.D a_27244_56974# 0.00166f
C529 xaa6.xe.XA1.MN0.G xaa6.xe.XA7.MN2.D 2.12e-19
C530 xaa6.xd.XA7.MP1.G a_29764_57326# 9.02e-20
C531 xaa6.xf.XA7.MN1.G xaa6.xf.XA7.MN0.D 0.0449f
C532 xaa6.xd.XA7.MN1.G a_28612_57326# 0.00174f
C533 xaa6.xc.XA1.MN0.G a_26092_56974# 1.06e-19
C534 AVDD a_31132_55918# 0.00151f
C535 xaa6.xc.XA5.MN0.G xaa6.xd.XA5.MN0.G 0.00217f
C536 xaa6.xe.XA7.MN1.D a_32284_53454# 6.39e-19
C537 xaa6.xe.XA1.MN0.G a_31132_53454# 0.0778f
C538 a_32284_55918# a_32284_55566# 0.0109f
C539 xaa1.xa4.M0.D m1_4468_100124# 67.7f
C540 xaa1.xa4.M0.D m3_4788_88764# 0.0138f
C541 xaa4.xa1.M4.D xaa4.xa1.M3.D 0.0488f
C542 a_36172_54158# a_36172_53806# 0.0109f
C543 a_4308_53678# xbb1.xa3.M7.D 0.00155f
C544 li_4468_97084# li_4468_96284# 39.3f
C545 a_n508_74698# xaa1.xa4.M0.D 3.69e-19
C546 a_27244_58030# xaa6.xc.XA7.MN1.D 0.0658f
C547 a_26092_58030# xaa6.xc.XA1.MN0.G 1.35e-19
C548 CK a_37324_56622# 8.7e-19
C549 xaa1.xa3.D a_10092_55566# 0.0702f
C550 AVDD a_244_56270# 0.384f
C551 xaa6.xf.XA7.MN1.G xaa6.xf.XA4.MN0.D 1.09e-19
C552 a_31132_56974# xaa6.xe.XA5.MN0.G 1.67e-19
C553 xaa6.xd.XA6.MP0.D a_28612_56270# 0.0467f
C554 xaa6.xf.XA1.MN0.G a_34804_54862# 0.00233f
C555 xaa6.xd.XA7.MP1.G a_28612_55214# 0.027f
C556 xaa6.xd.XA7.MN1.G a_27244_55214# 7.1e-20
C557 xaa6.xc.XA1.MN0.G xaa6.xd.XA3.MP0.D 0.00218f
C558 AVDD a_27244_53454# 0.367f
C559 a_36172_54862# a_36172_54510# 0.0109f
C560 xaa6.xd.XA3.MP0.D a_29764_54510# 2.16e-19
C561 xaa6.xd.XA3.MN0.D a_28612_54510# 2.16e-19
C562 xaa1.xa4.M0.D m3_37668_105244# 0.074f
C563 xaa4.xa2.M0.G m3_22620_58180# 0.0273f
C564 xaa1.xa4.M0.D a_n908_63622# 0.00697f
C565 a_1220_70022# a_2948_70022# 9.03e-19
C566 AVDD a_5844_58494# 0.348f
C567 CK xaa6.xg.XA7.MN1.D 0.00311f
C568 xaa0.xa6.MN0.D a_n908_56622# 0.00338f
C569 xaa5.xa3.xc1a.D a_27244_60750# 0.00176f
C570 m2_4468_107804# m3_37748_108124# 0.0138f
C571 a_n908_56622# xaa0.xa1.MN0.G 7.25e-20
C572 a_32284_56974# a_33652_56974# 8.89e-19
C573 xaa0.xa5.MN0.D a_n908_55918# 0.0799f
C574 xaa6.xe.XA1.MN0.G a_33652_55918# 0.00209f
C575 xaa6.xf.XA7.MN1.G xaa6.xf.XA6.MN0.D 0.0158f
C576 PWRUP_1V8 a_31132_54862# 0.00561f
C577 xaa6.xd.XA7.MN1.G a_29764_56270# 0.00344f
C578 xaa0.xa3.MN1.G a_n908_55566# 0.0895f
C579 AVDD a_33652_54862# 0.383f
C580 xaa1.xa4.M0.D m2_4468_86684# 71.5f
C581 AVDD li_6132_61812# 0.00142f
C582 a_27244_53102# a_28612_53102# 8.89e-19
C583 li_4468_79964# li_4468_79804# 7.91f
C584 xaa5.xb2_1.MN0.D xaa5.xb2_0.MN0.D 0.197f
C585 AVDD CK 3.95f
C586 a_36172_57678# a_36172_57326# 0.0109f
C587 xaa6.xc.XA7.MN1.D a_26092_56974# 0.0092f
C588 xaa0.xa5.MN2.G a_27244_56974# 0.0725f
C589 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MN2.D 0.0372f
C590 xaa6.xd.XA7.MP1.G a_28612_57326# 0.0948f
C591 xaa6.xf.XA7.MP1.G xaa6.xf.XA7.MN0.D 0.117f
C592 AVDD a_29764_55918# 0.00151f
C593 xaa6.xd.XA7.MN1.G a_29764_53806# 0.115f
C594 xaa6.xd.XA1.MN0.G a_32284_53454# 1.11e-19
C595 xaa4.xa2.M0.D xaa4.xa1.M8.D 0.206f
C596 xaa1.xa4.M0.D m1_4468_101084# 67.7f
C597 xaa1.xa4.M0.D m3_4628_88764# 0.0276f
C598 xaa3.xa1b.MN0.D xaa3.xa5a.MN0.D 0.224f
C599 IBPSR_1U xaa1.xa2.M3.D 0.026f
C600 a_356_74698# a_1220_74698# 0.071f
C601 m1_4468_109724# m2_4468_109724# 12.9f
C602 AVDD a_n908_56270# 0.00159f
C603 a_32284_58030# a_33652_58030# 8.89e-19
C604 a_27244_58030# xaa0.xa5.MN2.G 0.0337f
C605 a_26092_58030# xaa6.xc.XA7.MN1.D 0.0709f
C606 PWRUP_1V8 xaa0.xa5.MN0.D 0.00513f
C607 m2_4468_94364# m3_37748_94684# 0.0138f
C608 xaa6.xf.XA7.MP1.G xaa6.xf.XA4.MN0.D 0.056f
C609 xaa6.xf.XA7.MN1.G xaa6.xf.XA4.MP0.D 0.00941f
C610 PWRUP_1V8 xaa4.xa1.M1.D 9.97e-19
C611 xaa1.xa4.M0.D li_4468_89404# 23f
C612 xaa6.xf.XA6.MP0.D xaa6.xf.XA6.MN0.D 0.00918f
C613 xaa6.xf.XA7.MN1.D a_34804_54862# 0.00652f
C614 xaa6.xf.XA1.MN0.G a_33652_54862# 1.35e-19
C615 xaa6.xc.XA1.MN0.G xaa6.xc.XA3.MP0.D 0.00238f
C616 AVDD a_26092_53454# 0.00159f
C617 xaa6.xd.XA3.MP0.D a_28612_54510# 0.0467f
C618 xaa1.xa4.M0.D m3_4788_106044# 0.0138f
C619 a_37324_55566# m1_37504_55818# 0.0131f
C620 li_4468_114364# li_4468_113564# 39.3f
C621 xaa4.xa2.M0.G m3_22548_58180# 0.0137f
C622 a_1652_72222# xaa1.xa3.D 0.168f
C623 li_4468_80924# m1_4468_80924# 23f
C624 xaa1.xa1.M3.D xaa1.xa1.M2.D 0.0488f
C625 xaa0.xa6.MN0.D xaa0.xa3.MN1.G 0.142f
C626 CK xaa6.xf.XA1.MN0.G 0.0445f
C627 AVDD a_4692_58494# 0.00171f
C628 m2_4468_107804# m3_37668_108124# 0.0138f
C629 xaa0.xa5.MN0.D xaa0.xa5.MP1.D 0.0657f
C630 a_26092_56974# a_26092_56622# 0.0109f
C631 xaa6.xe.XA7.MN2.D a_31132_56622# 0.00176f
C632 xaa0.xa3.MN1.G xaa0.xa1.MN0.G 0.439f
C633 xaa6.xe.XA1.MN0.G a_32284_55918# 0.0022f
C634 xaa6.xf.XA7.MP1.G xaa6.xf.XA6.MN0.D 0.056f
C635 xaa6.xf.XA7.MN1.G xaa6.xf.XA6.MP0.D 0.0285f
C636 PWRUP_1V8 a_29764_54862# 0.00561f
C637 xaa6.xd.XA7.MP1.G a_29764_56270# 0.1f
C638 xaa6.xd.XA7.MN1.G a_28612_56270# 0.0803f
C639 AVDD a_32284_54862# 0.383f
C640 xaa1.xa4.M0.D m2_4468_87644# 71.5f
C641 xaa6.xc.XA4.MN0.D a_26092_55214# 0.0472f
C642 xaa6.xe.XA5.MN0.G xaa6.xe.XA3.MP0.D 0.0488f
C643 a_34804_53454# a_34804_53102# 0.0109f
C644 CK xaa5.xb1.MN1.D 7.29e-20
C645 xaa5.xa3.xb1_0.D xaa5.xb2_0.MN0.D 0.00359f
C646 xaa3.xa1b.MN0.D xaa3.xa3a.MN0.D 0.224f
C647 IBPSR_1U xaa1.xb1.M0.D 8.96e-19
C648 a_27244_62158# a_28612_62158# 8.89e-19
C649 xaa1.xa2.M2.D xaa1.xa2.M1.D 0.0488f
C650 AVDD a_29764_62862# 0.00139f
C651 m1_4468_76124# m2_4468_76124# 12.9f
C652 PWRUP_1V8 a_26092_55918# 0.00675f
C653 xaa0.xa5.MN2.G a_26092_56974# 0.066f
C654 xaa6.xf.XA7.MP1.G xaa6.xf.XA7.MN1.G 0.537f
C655 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN2.D 0.00981f
C656 AVDD a_28612_55918# 0.385f
C657 m2_4468_80924# m3_37748_81244# 0.0138f
C658 xaa6.xd.XA7.MN1.G a_28612_53806# 0.113f
C659 xaa6.xd.XA7.MP1.G a_29764_53806# 0.00375f
C660 xaa6.xd.XA1.MN0.G a_31132_53454# 0.00212f
C661 a_31132_55918# a_31132_55566# 0.0109f
C662 xaa1.xa4.M0.D m1_4468_102044# 67.7f
C663 xaa1.xa4.M0.D m3_37748_88924# 0.111f
C664 a_34804_54158# a_34804_53806# 0.0109f
C665 li_4468_97244# li_4468_97084# 7.91f
C666 xaa1.xa3.D xaa1.xa2.M2.D 0.00119f
C667 a_n908_63270# xaa1.xa2.M3.D 1.21e-19
C668 xbb0.xa1.XA1.N xaa1.xa4.M0.D 0.448f
C669 a_26092_58030# xaa0.xa5.MN2.G 0.0473f
C670 AVDD xaa0.xa5.MN2.D 0.00193f
C671 m2_4468_94364# m3_37668_94684# 0.0138f
C672 xaa6.xc.XA6.MP0.D a_27244_56270# 0.0467f
C673 a_29764_56974# xaa6.xd.XA5.MN0.G 1.55e-19
C674 xaa6.xf.XA7.MP1.G xaa6.xf.XA4.MP0.D 0.0615f
C675 xaa4.xa4.M0.D xaa4.xa1.M5.D 5.55e-19
C676 PWRUP_1V8 xaa6.xg.XA1.MN0.D 0.0103f
C677 xaa6.xc.XA7.MN1.D xaa6.xc.XA3.MP0.D 0.0844f
C678 xaa6.xf.XA7.MN1.D a_33652_54862# 0.00464f
C679 xaa6.xe.XA1.MN0.G a_34804_54862# 1.02e-19
C680 xaa6.xc.XA1.MN0.G xaa6.xc.XA3.MN0.D 6.01e-19
C681 a_34804_54862# a_34804_54510# 0.0109f
C682 xaa1.xa4.M0.D m3_4628_106044# 0.0276f
C683 PWRUP_1V8 m1_37504_55818# 3.46e-19
C684 xaa4.xa2.M0.G m3_13116_58356# 0.0634f
C685 a_1220_70022# xaa1.xa3.D 0.0035f
C686 a_4692_60782# a_5844_60782# 0.00133f
C687 PWRUP_1V8 a_n908_59750# 1.28e-19
C688 xaa0.xa6.MN0.D a_244_56974# 0.0313f
C689 CK xaa6.xf.XA7.MN1.D 2.93e-19
C690 AVDD a_11712_59086# 0.424f
C691 xaa0.xa3.MN1.G a_244_55918# 5.88e-19
C692 a_31132_56974# a_32284_56974# 0.00133f
C693 xaa6.xe.XA1.MN0.G a_31132_55918# 1.25e-19
C694 xaa6.xe.XA7.MN1.D a_32284_55918# 0.00149f
C695 xaa6.xf.XA7.MP1.G xaa6.xf.XA6.MP0.D 0.0619f
C696 AVDD a_31132_54862# 0.00151f
C697 xaa6.xd.XA7.MP1.G a_28612_56270# 0.0268f
C698 xaa6.xd.XA7.MN1.G a_27244_56270# 7.1e-20
C699 CK a_36172_54510# 2.59e-20
C700 xaa0.xa5.MN2.G xaa4.xa2.M0.D 7.16e-20
C701 xaa1.xa4.M0.D m2_4468_88604# 71.5f
C702 xaa6.xe.XA5.MN0.G xaa6.xe.XA3.MN0.D 0.0488f
C703 xaa1.xa4.M0.D m3_4788_72444# 0.0138f
C704 a_26092_53102# a_27244_53102# 0.00133f
C705 li_4468_103964# m1_4468_103964# 23f
C706 li_4468_80764# li_4468_79964# 39.3f
C707 xaa5.xa3.xb1_0.D xaa5.xa3.xc2a.D 0.0467f
C708 IBPSR_1U xaa3.xa3a.MN0.D 3.69e-20
C709 AVDD a_28612_62862# 0.352f
C710 xaa4.xa2.M0.G a_10092_55038# 0.0708f
C711 a_34804_57678# a_34804_57326# 0.0109f
C712 xaa6.xc.XA7.MN0.D a_27244_57326# 0.0525f
C713 AVDD a_27244_55918# 0.385f
C714 m2_4468_80924# m3_37668_81244# 0.0138f
C715 xaa6.xd.XA1.MN0.G a_29764_53454# 0.0733f
C716 xaa6.xd.XA7.MN1.G a_27244_53806# 7.1e-20
C717 xaa6.xd.XA7.MP1.G a_28612_53806# 0.00282f
C718 a_37324_55918# xaa6.xg.XA5.MN0.G 0.0658f
C719 xaa1.xa4.M0.D m1_4468_103004# 67.7f
C720 xaa1.xa4.M0.D m3_37668_88924# 0.074f
C721 IBPSR_1U xaa1.xa2.M4.D 0.026f
C722 a_29764_63566# xaa5.xb2_4.MN0.D 0.0682f
C723 a_n940_74698# xaa1.xa4.M0.D 0.187f
C724 m1_4468_110684# m2_4468_110684# 12.9f
C725 a_31132_58030# a_32284_58030# 0.00133f
C726 PWRUP_1V8 a_n908_56622# 7.32e-19
C727 AVDD xaa0.xa5.MN0.D 0.697f
C728 xaa6.xc.XA6.MP0.D a_26092_56270# 2.16e-19
C729 xaa6.xc.XA6.MN0.D a_27244_56270# 2.16e-19
C730 xaa6.xc.XA7.MP1.G a_27244_55214# 0.027f
C731 xaa6.xc.XA7.MN1.G a_28612_55214# 7.1e-20
C732 xaa4.xa4.M0.D xaa4.xa1.M6.D 5.76e-19
C733 PWRUP_1V8 xaa6.xf.XA1.MN0.D 0.0103f
C734 xaa1.xa4.M0.D li_4468_90364# 23f
C735 xaa6.xc.XA7.MN1.D xaa6.xc.XA3.MN0.D 0.0425f
C736 xaa6.xe.XA1.MN0.G a_33652_54862# 0.00209f
C737 AVDD xaa4.xa1.M1.D 0.00415f
C738 xaa6.xg.XA7.MN0.G xaa6.xg.XA5.MN0.G 9.76e-20
C739 xaa6.xc.XA3.MP0.D a_27244_54510# 0.0467f
C740 xaa6.xf.XA3.MP0.D xaa6.xf.XA3.MN0.D 0.00918f
C741 xaa1.xa4.M0.D m3_37748_106204# 0.111f
C742 PWRUP_1V8 m1_37504_57930# 0.00289f
C743 li_4468_114524# li_4468_114364# 7.91f
C744 xaa4.xa2.M0.G m3_13044_58356# 0.106f
C745 a_1220_70022# a_2084_70022# 0.071f
C746 a_788_72222# a_2948_70022# 2.35e-20
C747 a_640_60806# xaa1.xb2.M0.D 0.00155f
C748 PWRUP_1V8 xaa4.xa4.M0.D 0.00178f
C749 xaa1.xa1.M7.D a_n908_59750# 5.02e-20
C750 xaa1.xa1.M8.D a_640_59750# 0.0729f
C751 xaa0.xa6.MN0.D a_n908_56974# 0.0312f
C752 CK xaa6.xe.XA1.MN0.G 0.064f
C753 xaa0.xa2a.MN0.D xaa1.xa1.M0.D 0.00139f
C754 AVDD a_640_59750# 0.389f
C755 xaa6.xd.XA1.MN0.G a_32284_55918# 1.11e-19
C756 xaa6.xd.XA7.MN2.D a_29764_56622# 0.00176f
C757 xaa0.xa3.MN1.G a_n908_55918# 0.0367f
C758 xaa6.xe.XA7.MN1.D a_31132_55918# 0.00829f
C759 AVDD a_29764_54862# 0.00151f
C760 xaa1.xa4.M0.D m2_4468_89564# 71.5f
C761 xaa4.xa1.M8.D a_10092_54510# 0.0541f
C762 a_11712_55918# a_11712_54334# 0.00223f
C763 xaa1.xa4.M0.D m3_4628_72444# 0.0276f
C764 a_37324_56622# m1_37504_55818# 5.6e-19
C765 a_33652_53454# a_33652_53102# 0.0109f
C766 xaa5.xb2_1.MN0.D a_29764_62158# 0.126f
C767 IBPSR_1U xaa1.xa1.M0.D 0.0288f
C768 a_26092_62158# a_27244_62158# 0.00133f
C769 AVDD a_27244_62862# 0.469f
C770 m1_4468_77084# m2_4468_77084# 12.9f
C771 xaa6.xc.XA7.MN0.D a_26092_57326# 0.055f
C772 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MN2.D 0.0372f
C773 PWRUP_1V8 xaa6.xg.XA6.MN0.G 0.0294f
C774 xaa6.xe.XA7.MP1.G xaa6.xf.XA7.MN1.G 1.74e-19
C775 xaa6.xc.XA7.MP1.G a_27244_57326# 0.0964f
C776 AVDD a_26092_55918# 0.00159f
C777 xaa6.xd.XA1.MN0.G a_28612_53454# 0.0676f
C778 a_37324_55918# xaa6.xg.XA5.MN0.D 0.0215f
C779 a_36172_55918# xaa6.xg.XA5.MN0.G 0.0731f
C780 a_29764_55918# a_29764_55566# 0.0109f
C781 xaa1.xa4.M0.D m1_4468_103964# 67.7f
C782 xaa6.xg.XA7.MN1.D m1_37504_55818# 0.0772f
C783 xaa1.xa4.M0.D m3_4788_89724# 0.0138f
C784 a_33652_54158# a_33652_53806# 0.0109f
C785 li_4468_98044# li_4468_97244# 39.3f
C786 a_n908_63270# xaa1.xa2.M4.D 1.81e-19
C787 a_28612_63566# xaa5.xb2_4.MN0.D 0.0674f
C788 xaa3.xa1b.MN0.D a_4692_62718# 0.00468f
C789 AVDD xaa1.xa4.M0.D 0.873f
C790 PWRUP_1V8 xaa0.xa3.MN1.G 0.0502f
C791 AVDD a_244_56622# 0.388f
C792 xaa6.xc.XA6.MN0.D a_26092_56270# 0.0474f
C793 xaa6.xc.XA7.MP1.G a_26092_55214# 0.0944f
C794 xaa6.xc.XA7.MN1.G a_27244_55214# 0.0761f
C795 xaa4.xa4.M0.D a_11712_54334# 0.0198f
C796 PWRUP_1V8 xaa6.xe.XA1.MN0.D 0.0103f
C797 xaa6.xe.XA1.MN0.G a_32284_54862# 0.00257f
C798 AVDD xaa6.xg.XA1.MN0.D 2.4e-19
C799 a_33652_54862# a_33652_54510# 0.0109f
C800 xaa6.xc.XA3.MN0.D a_27244_54510# 2.16e-19
C801 xaa6.xc.XA3.MP0.D a_26092_54510# 2.16e-19
C802 xaa1.xa4.M0.D m3_37668_106204# 0.074f
C803 AVDD m1_37504_55818# 0.427f
C804 xaa4.xa2.M0.G m3_22620_59236# 0.0273f
C805 li_4468_81884# m1_4468_81884# 23f
C806 CK xaa6.xe.XA7.MN1.D 9.13e-19
C807 xaa0.xa2a.MN0.D a_640_60278# 6.01e-19
C808 AVDD a_n908_59750# 0.00649f
C809 xaa6.xd.XA1.MN0.G a_31132_55918# 0.00205f
C810 xaa0.xa3.MN1.G xaa0.xa5.MP1.D 0.00164f
C811 xaa6.xg.XA7.MN0.G a_37324_56974# 0.0674f
C812 a_29764_56974# a_31132_56974# 8.89e-19
C813 xaa6.xg.XA7.MN2.D a_36172_56974# 0.0494f
C814 PWRUP_1V8 a_26092_54862# 0.00554f
C815 AVDD a_28612_54862# 0.383f
C816 xaa1.xa4.M0.D m2_4468_90524# 71.5f
C817 xaa6.xd.XA5.MN0.G xaa6.xd.XA3.MN0.D 0.0488f
C818 xaa1.xa4.M0.D m3_37748_72604# 0.111f
C819 a_37324_56622# m1_37504_57930# 8.83e-19
C820 li_4468_80924# li_4468_80764# 7.91f
C821 CK a_29764_61806# 3.97e-20
C822 xaa5.xb2_1.MN0.D a_28612_62158# 0.0878f
C823 IBPSR_1U a_640_60278# 0.00122f
C824 AVDD a_26092_62862# 0.00168f
C825 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN2.D 0.0101f
C826 PWRUP_1V8 xaa6.xf.XA6.MN0.G 0.0466f
C827 xaa6.xe.XA7.MN1.G xaa6.xf.XA7.MN1.G 0.31f
C828 xaa6.xe.XA7.MP1.G xaa6.xf.XA7.MP1.G 0.00435f
C829 a_33652_57678# a_33652_57326# 0.0109f
C830 xaa6.xc.XA7.MP1.G a_26092_57326# 9.02e-20
C831 xaa6.xc.XA7.MN1.G a_27244_57326# 0.00174f
C832 AVDD a_11712_55918# 0.424f
C833 xaa6.xc.XA1.MN0.G a_29764_53454# 1.02e-19
C834 xaa6.xd.XA7.MN1.D a_28612_53454# 6.39e-19
C835 a_36172_55918# xaa6.xg.XA5.MN0.D 0.0215f
C836 xaa1.xa4.M0.D m1_4468_104924# 67.7f
C837 xaa6.xf.XA1.MN0.G xaa6.xg.XA1.MN0.D 0.00287f
C838 xaa6.xg.XA7.MN1.D m1_37504_57930# 0.0757f
C839 xaa1.xa4.M0.D m3_4628_89724# 0.0276f
C840 xaa6.xg.XA3.MN1.G a_37324_53454# 0.0767f
C841 a_37324_54510# m1_37504_55818# 8.83e-19
C842 a_29764_64270# CK 7.76e-19
C843 xaa5.xa3.xb2_0.G xaa5.xb2_4.MN0.D 0.228f
C844 a_28612_63566# a_29764_63566# 0.00133f
C845 m1_4468_111644# m2_4468_111644# 12.9f
C846 a_29764_58030# a_31132_58030# 8.89e-19
C847 xaa1.xa3.D xaa4.xa2.M0.D 0.00551f
C848 AVDD a_n908_56622# 0.00171f
C849 xaa6.xe.XA6.MN0.D xaa6.xe.XA6.MP0.D 0.00918f
C850 xaa6.xc.XA7.MN1.G a_26092_55214# 0.00134f
C851 xaa4.xa4.M0.D xaa4.xa1.M7.D 6.08e-19
C852 PWRUP_1V8 xaa6.xd.XA1.MN0.D 0.0103f
C853 xaa1.xa4.M0.D li_4468_91324# 23f
C854 xaa6.xe.XA7.MN1.D a_32284_54862# 0.00464f
C855 xaa6.xe.XA1.MN0.G a_31132_54862# 4.77e-19
C856 xaa6.xe.XA7.MP1.G xaa6.xe.XA4.MP0.D 0.0615f
C857 AVDD xaa6.xf.XA1.MN0.D 2.4e-19
C858 AVDD m1_37504_57930# 0.329f
C859 xaa6.xc.XA3.MN0.D a_26092_54510# 0.0474f
C860 xaa1.xa4.M0.D m3_4788_107004# 0.0138f
C861 li_4468_115324# li_4468_114524# 39.3f
C862 xaa4.xa2.M0.G m3_22548_59236# 0.0137f
C863 a_788_72222# xaa1.xa3.D 0.0413f
C864 xaa1.xb2.M7.D xaa1.xb2.M0.D 0.0488f
C865 CK xaa6.xd.XA1.MN0.G 8.66e-19
C866 PWRUP_1V8 a_29764_60750# 0.078f
C867 xaa0.xa2a.MN0.D xaa1.xa1.M1.D 0.0019f
C868 AVDD xaa4.xa4.M0.D 11.4f
C869 m2_4468_108764# m3_37748_109084# 0.0138f
C870 xaa6.xc.XA7.MP1.G a_27244_56270# 0.0268f
C871 xaa6.xc.XA7.MN1.G a_28612_56270# 7.1e-20
C872 xaa6.xg.XA7.MN1.D xaa6.xg.XA6.MN0.G 0.027f
C873 xaa6.xd.XA1.MN0.G a_29764_55918# 0.00217f
C874 xaa6.xg.XA7.MN0.G a_36172_56974# 0.0658f
C875 PWRUP_1V8 xaa6.xg.XA4.MN0.G 0.0154f
C876 xaa6.xe.XA7.MP1.G xaa6.xe.XA6.MP0.D 0.0619f
C877 AVDD a_27244_54862# 0.383f
C878 xaa6.xd.XA5.MN0.G xaa6.xd.XA3.MP0.D 0.0488f
C879 xaa1.xa4.M0.D m2_4468_91484# 71.5f
C880 xaa6.xg.XA5.MN0.G a_37324_54862# 0.0225f
C881 a_37324_55566# a_37324_55214# 0.0109f
C882 xaa1.xa4.M0.D m3_37668_72604# 0.074f
C883 a_32284_53454# a_32284_53102# 0.0109f
C884 li_4468_104924# m1_4468_104924# 23f
C885 IBPSR_1U xaa1.xa1.M1.D 0.0267f
C886 xaa5.xa3.xb2_0.D a_27244_61806# 0.0303f
C887 AVDD xaa5.xb2_3.MN0.D 0.545f
C888 m1_4468_78044# m2_4468_78044# 12.9f
C889 xaa6.xc.XA1.MN0.G xaa6.xc.XA7.MN2.D 2.12e-19
C890 PWRUP_1V8 xaa6.xe.XA6.MN0.G 0.0465f
C891 xaa6.xe.XA7.MN1.G xaa6.xf.XA7.MP1.G 1.74e-19
C892 xaa6.xc.XA7.MN1.G a_26092_57326# 0.0781f
C893 xaa6.xe.XA7.MP1.G xaa6.xe.XA7.MN0.D 0.117f
C894 AVDD xaa6.xg.XA6.MN0.G 0.478f
C895 xaa6.xc.XA1.MN0.G a_28612_53454# 0.00209f
C896 a_4692_55150# a_5844_55150# 0.00133f
C897 xaa6.xf.XA6.MN0.G a_34804_55566# 0.00224f
C898 a_28612_55918# a_28612_55566# 0.0109f
C899 xaa1.xa4.M0.D m1_4468_105884# 67.7f
C900 xaa6.xc.XA7.MN1.G a_28612_53806# 7.1e-20
C901 xaa6.xc.XA7.MP1.G a_27244_53806# 0.00282f
C902 xaa6.xf.XA1.MN0.G xaa6.xf.XA1.MN0.D 0.0147f
C903 xaa1.xa4.M0.D m3_37748_89884# 0.111f
C904 xaa6.xf.XA1.MN0.G m1_37504_57930# 0.051f
C905 xaa6.xg.XA3.MN1.G a_36172_53454# 0.0148f
C906 a_n908_52750# a_244_52750# 0.00133f
C907 a_32284_54158# a_32284_53806# 0.0109f
C908 li_4468_98204# li_4468_98044# 7.91f
C909 xaa3.xa7.MN0.D a_4692_62366# 2.18e-19
C910 a_28612_64270# CK 0.00102f
C911 xaa3.xa1b.MN0.D xaa3.xa6.MN0.D 0.137f
C912 xaa5.xa3.xb2_0.G a_29764_63566# 0.134f
C913 IBPSR_1U xaa1.xa2.M5.D 0.026f
C914 PWRUP_1V8 a_n908_56974# 8.53e-19
C915 AVDD xaa0.xa3.MN1.G 1.25f
C916 m2_4468_95324# m3_37748_95644# 0.0138f
C917 a_26092_56974# xaa6.xc.XA5.MN0.G 1.67e-19
C918 PWRUP_1V8 xaa6.xc.XA1.MN0.D 0.0107f
C919 CK a_37324_53102# 0.0692f
C920 xaa6.xe.XA7.MN1.D a_31132_54862# 0.00652f
C921 xaa6.xd.XA1.MN0.G a_32284_54862# 1.11e-19
C922 xaa6.xe.XA7.MP1.G xaa6.xe.XA4.MN0.D 0.056f
C923 xaa6.xe.XA7.MN1.G xaa6.xe.XA4.MP0.D 0.00941f
C924 AVDD xaa6.xe.XA1.MN0.D 1.75e-19
C925 a_32284_54862# a_32284_54510# 0.0109f
C926 xaa1.xa4.M0.D m3_4628_107004# 0.0276f
C927 xaa4.xa2.M0.G m3_13116_59412# 0.0634f
C928 xaa1.xa4.M0.D xaa1.xa4.M0.G 0.231f
C929 PWRUP_1V8 a_28612_60750# 0.0661f
C930 AVDD a_11712_60670# 0.362f
C931 m2_4468_108764# m3_37668_109084# 0.0138f
C932 xaa6.xd.XA1.MN0.G a_28612_55918# 1.35e-19
C933 xaa6.xc.XA7.MP1.G a_26092_56270# 0.0985f
C934 xaa6.xc.XA7.MN1.G a_27244_56270# 0.0819f
C935 xaa6.xd.XA7.MN1.D a_29764_55918# 0.00829f
C936 a_28612_56974# a_29764_56974# 0.00133f
C937 xaa6.xf.XA1.MN0.G xaa6.xg.XA6.MN0.G 0.00415f
C938 xaa6.xe.XA7.MP1.G xaa6.xe.XA6.MN0.D 0.056f
C939 xaa6.xe.XA7.MN1.G xaa6.xe.XA6.MP0.D 0.0285f
C940 AVDD a_26092_54862# 0.00159f
C941 xaa6.xg.XA5.MN0.G a_36172_54862# 0.033f
C942 xaa1.xa4.M0.D m2_4468_92444# 71.5f
C943 xaa4.xa1.M1.D a_10092_52750# 5.84e-19
C944 xaa1.xa4.M0.D m3_4788_73404# 0.0138f
C945 li_4468_81724# li_4468_80924# 39.3f
C946 xaa5.xa3.xb1_0.D a_27244_62158# 0.14f
C947 a_29764_62510# a_29764_62158# 0.0109f
C948 xaa3.xa1b.MN0.D a_4692_60430# 0.00455f
C949 xaa5.xa3.xb2_0.D a_26092_61806# 0.0351f
C950 AVDD a_29764_63214# 0.00139f
C951 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MN2.D 0.0372f
C952 PWRUP_1V8 xaa6.xd.XA6.MN0.G 0.0466f
C953 a_32284_57678# a_32284_57326# 0.0109f
C954 xaa6.xe.XA7.MN1.G xaa6.xe.XA7.MN0.D 0.0449f
C955 AVDD xaa6.xf.XA6.MN0.G 1.7f
C956 m2_4468_81884# m3_37748_82204# 0.0138f
C957 xaa6.xc.XA1.MN0.G a_27244_53454# 0.0739f
C958 a_34804_55918# xaa6.xf.XA5.MN0.G 0.0715f
C959 a_5844_55502# a_5844_55150# 0.0109f
C960 xaa6.xf.XA6.MN0.G a_33652_55566# 0.0154f
C961 xaa1.xa4.M0.D m1_4468_106844# 67.7f
C962 xaa6.xc.XA7.MP1.G a_26092_53806# 0.00375f
C963 xaa6.xc.XA7.MN1.G a_27244_53806# 0.115f
C964 xaa6.xg.XA7.MP1.G a_37324_54158# 0.0545f
C965 a_244_53102# a_244_52750# 0.0109f
C966 xaa1.xa4.M0.D m3_37668_89884# 0.074f
C967 xaa5.xa3.xb2_0.G a_28612_63566# 0.0958f
C968 xaa5.xb3.MP1.D CK 0.00519f
C969 a_n908_63270# xaa1.xa2.M5.D 2.99e-19
C970 a_29764_63918# a_29764_63566# 0.0109f
C971 m1_4468_112604# m2_4468_112604# 12.9f
C972 a_28612_58030# a_29764_58030# 0.00133f
C973 AVDD a_244_56974# 0.349f
C974 m2_4468_95324# m3_37668_95644# 0.0138f
C975 xaa6.xg.XA7.MN1.D xaa6.xg.XA4.MN0.G 0.028f
C976 CK a_36172_53102# 0.0761f
C977 xaa6.xd.XA1.MN0.G a_31132_54862# 0.00205f
C978 xaa6.xe.XA7.MN1.G xaa6.xe.XA4.MN0.D 1.09e-19
C979 xaa1.xa4.M0.D li_4468_92284# 23f
C980 AVDD xaa6.xd.XA1.MN0.D 2.4e-19
C981 xaa6.xe.XA3.MN0.D xaa6.xe.XA3.MP0.D 0.00918f
C982 xaa1.xa4.M0.D m3_37748_107164# 0.111f
C983 xaa4.xa2.M0.G m3_13044_59412# 0.106f
C984 li_4468_115484# li_4468_115324# 7.91f
C985 xaa1.xa4.M0.D a_n908_64150# 0.00719f
C986 li_4468_82844# m1_4468_82844# 23f
C987 xaa1.xa1.M4.D xaa1.xa1.M3.D 0.0488f
C988 AVDD a_29764_60750# 0.00511f
C989 xaa6.xc.XA1.MN0.G a_29764_55918# 1.02e-19
C990 xaa6.xc.XA7.MN1.G a_26092_56270# 0.00344f
C991 xaa6.xd.XA7.MN1.D a_28612_55918# 0.00149f
C992 xaa6.xf.XA7.MN2.D a_34804_56974# 0.0494f
C993 xaa6.xc.XA7.MN2.D a_26092_56622# 0.00176f
C994 PWRUP_1V8 a_36172_55214# 0.00579f
C995 xaa6.xf.XA1.MN0.G xaa6.xf.XA6.MN0.G 0.0112f
C996 xaa6.xe.XA7.MN1.G xaa6.xe.XA6.MN0.D 0.0158f
C997 AVDD xaa6.xg.XA4.MN0.G 0.485f
C998 xaa6.xc.XA5.MN0.G xaa6.xc.XA3.MP0.D 0.0488f
C999 a_36172_55566# a_36172_55214# 0.0109f
C1000 xaa1.xa4.M0.D m2_4468_93404# 71.5f
C1001 a_31132_53454# a_31132_53102# 0.0109f
C1002 xaa1.xa4.M0.D m3_4628_73404# 0.0276f
C1003 xaa5.xa4.MN0.D a_27244_62158# 0.00224f
C1004 xaa5.xa3.xb1_0.D a_26092_62158# 0.0809f
C1005 xaa3.xa1b.MN0.D xaa3.xa4.MN0.D 0.0558f
C1006 CK a_26092_61806# 1.18e-19
C1007 AVDD a_28612_63214# 0.352f
C1008 m1_4468_79004# m2_4468_79004# 12.9f
C1009 xaa0.xa5.MN2.G xaa6.xc.XA7.MN2.D 0.00981f
C1010 xaa6.xe.XA7.MN1.G xaa6.xe.XA7.MP1.G 0.537f
C1011 PWRUP_1V8 xaa6.xc.XA6.MN0.G 0.0462f
C1012 AVDD xaa6.xe.XA6.MN0.G 1.7f
C1013 m2_4468_81884# m3_37668_82204# 0.0138f
C1014 xaa6.xc.XA1.MN0.G a_26092_53454# 0.0778f
C1015 a_33652_55918# xaa6.xf.XA5.MN0.G 0.0674f
C1016 a_27244_55918# a_27244_55566# 0.0109f
C1017 xaa1.xa4.M0.D m1_4468_107804# 67.7f
C1018 xaa4.xa4.M0.D a_11712_52750# 0.00511f
C1019 xaa6.xc.XA7.MN1.G a_26092_53806# 0.114f
C1020 xaa4.xa2.M0.D a_10092_55566# 0.00102f
C1021 xaa6.xc.XA7.MN1.D a_27244_53454# 6.39e-19
C1022 xaa6.xe.XA1.MN0.G xaa6.xf.XA1.MN0.D 2.73e-19
C1023 xaa6.xg.XA7.MN1.G a_37324_54158# 0.0064f
C1024 xaa6.xg.XA7.MP1.G a_36172_54158# 0.057f
C1025 a_31132_54158# a_31132_53806# 0.0109f
C1026 xaa1.xa4.M0.D m3_4788_90684# 0.0138f
C1027 li_4468_99004# li_4468_98204# 39.3f
C1028 xaa0.xa6.MN0.D xaa1.xa2.M3.D 8.17e-19
C1029 xaa3.xa7.MN0.D xaa3.xa5a.MN0.D 0.00113f
C1030 a_29764_64622# CK 0.00192f
C1031 xaa3.xa1b.MN0.D a_5844_63070# 0.0677f
C1032 xaa4.xa2.M0.G xaa5.xb2_4.MN0.D 0.173f
C1033 IBPSR_1U xaa1.xa2.M6.D 0.026f
C1034 PWRUP_1V8 a_36172_57326# 0.00561f
C1035 AVDD a_n908_56974# 0.00623f
C1036 xaa6.xg.XA7.MN1.D a_37324_55214# 0.00145f
C1037 PWRUP_1V8 xaa4.xa1.M2.D 7.79e-19
C1038 CK a_34804_53102# 0.00126f
C1039 xaa6.xf.XA1.MN0.G xaa6.xg.XA4.MN0.G 0.00415f
C1040 xaa6.xd.XA1.MN0.G a_29764_54862# 0.00233f
C1041 AVDD xaa6.xc.XA1.MN0.D 1.75e-19
C1042 a_37324_54862# xaa6.xg.XA3.MP0.D 0.00176f
C1043 a_31132_54862# a_31132_54510# 0.0109f
C1044 xaa1.xa4.M0.D m3_37668_107164# 0.074f
C1045 xaa4.xa2.M0.G m3_22620_60292# 0.0273f
C1046 xaa5.xb1.MN1.D a_29764_60750# 4.81e-19
C1047 AVDD a_28612_60750# 0.336f
C1048 xaa6.xc.XA1.MN0.G a_28612_55918# 0.00209f
C1049 a_27244_56974# a_28612_56974# 8.89e-19
C1050 xaa3.xa1b.MN0.D xbb1.xa3.M7.D 1.38e-19
C1051 PWRUP_1V8 a_34804_55214# 0.00579f
C1052 xaa6.xf.XA7.MN1.D xaa6.xf.XA6.MN0.G 0.224f
C1053 AVDD a_37324_55214# 0.364f
C1054 xaa6.xc.XA5.MN0.G xaa6.xc.XA3.MN0.D 0.0488f
C1055 xaa1.xa4.M0.D m2_4468_94364# 71.5f
C1056 xaa1.xa4.M0.D m3_37748_73564# 0.111f
C1057 li_4468_81884# li_4468_81724# 7.91f
C1058 li_4468_105884# m1_4468_105884# 23f
C1059 xaa5.xa4.MN0.D a_26092_62158# 0.00224f
C1060 a_28612_62510# a_28612_62158# 0.0109f
C1061 AVDD a_27244_63214# 0.439f
C1062 xaa0.xa5.MN2.G a_244_56270# 0.0658f
C1063 xaa6.xg.XA7.MN1.D a_37324_57326# 0.00337f
C1064 a_37324_57678# xaa6.xg.XA7.MN0.D 0.00176f
C1065 a_31132_57678# a_31132_57326# 0.0109f
C1066 AVDD xaa6.xd.XA6.MN0.G 1.7f
C1067 xaa6.xe.XA6.MN0.G a_32284_55566# 0.0154f
C1068 xaa1.xa4.M0.D m1_4468_108764# 67.7f
C1069 a_4692_55502# a_4692_55150# 0.0109f
C1070 xaa6.xe.XA1.MN0.G xaa6.xe.XA1.MN0.D 0.0357f
C1071 xaa6.xg.XA7.MN1.G a_36172_54158# 2.31e-19
C1072 a_n908_53102# a_n908_52750# 0.0109f
C1073 xaa1.xa4.M0.D m3_4628_90684# 0.0276f
C1074 a_29764_63918# xaa5.xa3.xb2_0.G 0.0683f
C1075 a_28612_63918# a_28612_63566# 0.0109f
C1076 a_28612_64622# CK 0.00188f
C1077 xaa5.xb3.MP1.D a_28612_62862# 6e-20
C1078 a_n908_63270# xaa1.xa2.M6.D 5.84e-19
C1079 xaa3.xa1b.MN0.D a_4692_63070# 0.0743f
C1080 xaa4.xa2.M0.G a_29764_63566# 3.48e-19
C1081 m1_4468_113564# m2_4468_113564# 12.9f
C1082 PWRUP_1V8 a_34804_57326# 0.00567f
C1083 a_27244_58030# a_28612_58030# 8.89e-19
C1084 AVDD a_37324_57326# 0.364f
C1085 xaa6.xd.XA6.MP0.D xaa6.xd.XA6.MN0.D 0.00918f
C1086 xaa6.xg.XA7.MN1.D a_36172_55214# 0.00558f
C1087 PWRUP_1V8 a_37324_53806# 0.0658f
C1088 a_33652_56622# xaa6.xf.XA6.MN0.G 5.6e-19
C1089 xaa6.xf.XA1.MN0.G a_37324_55214# 1.11e-19
C1090 xaa6.xd.XA7.MN1.D a_29764_54862# 0.00652f
C1091 xaa6.xd.XA1.MN0.G a_28612_54862# 1.35e-19
C1092 xaa1.xa4.M0.D li_4468_93244# 23f
C1093 xaa1.xa4.M0.D m3_4788_107964# 0.0138f
C1094 xaa4.xa2.M0.G m3_22548_60292# 0.0137f
C1095 li_4468_116284# li_4468_115484# 39.3f
C1096 a_788_72222# a_1652_72222# 0.107f
C1097 a_n76_72222# xaa1.xa3.D 0.0376f
C1098 xaa1.xb2.M7.D a_640_60806# 0.0534f
C1099 xaa5.xb1.MN1.D a_28612_60750# 0.00224f
C1100 xaa0.xa2a.MN0.D xaa1.xa1.M2.D 0.0027f
C1101 AVDD a_27244_60750# 0.367f
C1102 xaa6.xc.XA1.MN0.G a_27244_55918# 0.0022f
C1103 IBPSR_1U xbb1.xa3.M7.D 0.0974f
C1104 xaa6.xe.XA1.MN0.G xaa6.xf.XA6.MN0.G 0.0181f
C1105 AVDD a_36172_55214# 0.00151f
C1106 xaa6.xf.XA5.MN0.G a_34804_54862# 0.033f
C1107 a_34804_55566# a_34804_55214# 0.0109f
C1108 xaa1.xa4.M0.D m2_4468_95324# 71.5f
C1109 xbb1.xa3.M7.D a_4308_51918# 5.02e-20
C1110 a_29764_53454# a_29764_53102# 0.0109f
C1111 xaa1.xa4.M0.D m3_37668_73564# 0.074f
C1112 IBPSR_1U xaa1.xa1.M2.D 0.0264f
C1113 xaa5.xa3.xb1_0.D xaa5.xb2_1.MN0.D 0.00229f
C1114 CK xaa5.xb2_0.MN0.D 7.29e-20
C1115 xaa5.xa3.xb2_0.D xaa5.xa3.xc2a.D 0.123f
C1116 AVDD a_26092_63214# 0.00154f
C1117 m1_4468_79964# m2_4468_79964# 12.9f
C1118 xaa0.xa5.MN2.G a_n908_56270# 0.0725f
C1119 a_37324_57678# xaa6.xg.XA7.MP1.G 0.0694f
C1120 PWRUP_1V8 a_36172_56270# 0.00783f
C1121 xaa6.xg.XA7.MN1.D a_36172_57326# 0.014f
C1122 a_36172_57678# xaa6.xg.XA7.MN0.D 0.00176f
C1123 AVDD xaa6.xc.XA6.MN0.G 1.7f
C1124 xaa6.xe.XA6.MN0.G a_31132_55566# 0.00224f
C1125 a_26092_55918# a_26092_55566# 0.0109f
C1126 xaa1.xa4.M0.D m1_4468_109724# 67.7f
C1127 a_4692_55502# a_5844_55502# 0.00133f
C1128 a_32284_55918# xaa6.xe.XA5.MN0.G 0.0658f
C1129 a_n908_53102# a_244_53102# 0.00133f
C1130 a_29764_54158# a_29764_53806# 0.0109f
C1131 xaa1.xa4.M0.D m3_37748_90844# 0.111f
C1132 li_4468_99164# li_4468_99004# 7.91f
C1133 xaa0.xa6.MN0.D xaa1.xa2.M4.D 8.17e-19
C1134 xaa3.xa7.MN0.D a_5844_62718# 0.00224f
C1135 xaa4.xa2.M0.G a_28612_63566# 0.0346f
C1136 a_28612_63918# xaa5.xa3.xb2_0.G 0.0674f
C1137 xaa5.xa3.xb1_0.G a_29764_63566# 0.00356f
C1138 xaa5.xb1.MN1.G xaa5.xb2_4.MN0.D 0.0401f
C1139 a_4692_63422# xaa3.xa6.MN0.D 7.11e-19
C1140 CK a_37324_56974# 8.62e-19
C1141 AVDD a_36172_57326# 0.00151f
C1142 xaa6.xf.XA1.MN0.G a_36172_55214# 0.00193f
C1143 a_37324_56622# a_37324_56270# 0.0109f
C1144 xaa6.xd.XA7.MN1.G xaa6.xd.XA4.MN0.D 1.09e-19
C1145 xaa6.xd.XA7.MN1.D a_28612_54862# 0.00464f
C1146 xaa6.xc.XA1.MN0.G a_29764_54862# 1.02e-19
C1147 PWRUP_1V8 a_36172_53806# 0.0753f
C1148 AVDD xaa4.xa1.M2.D 0.00415f
C1149 xaa4.xa2.M0.D xaa4.xa1.M0.D 8.24e-19
C1150 a_36172_54862# xaa6.xg.XA3.MN0.D 0.00176f
C1151 a_29764_54862# a_29764_54510# 0.0109f
C1152 xaa1.xa4.M0.D m3_4628_107964# 0.0276f
C1153 a_4692_57790# li_4980_56708# 4.95e-20
C1154 xaa4.xa2.M0.G m3_13116_60468# 0.0634f
C1155 li_4468_83804# m1_4468_83804# 23f
C1156 CK a_37324_58030# 0.00188f
C1157 AVDD a_26092_60750# 0.00543f
C1158 m2_4468_109724# m3_37748_110044# 0.0138f
C1159 xaa6.xc.XA1.MN0.G a_26092_55918# 1.25e-19
C1160 xaa6.xg.XA7.MN1.D a_37324_56270# 0.00378f
C1161 a_26092_56974# a_27244_56974# 0.00133f
C1162 IBPSR_1U xaa4.xa1.M3.D 0.026f
C1163 xaa6.xe.XA1.MN0.G xaa6.xe.XA6.MN0.G 0.0125f
C1164 xaa6.xd.XA7.MN1.G xaa6.xd.XA6.MN0.D 0.0158f
C1165 xaa6.xc.XA7.MN1.D a_27244_55918# 0.00149f
C1166 AVDD a_34804_55214# 0.00151f
C1167 xaa6.xf.XA6.MN0.G a_33652_54510# 0.00119f
C1168 xaa6.xf.XA5.MN0.G a_33652_54862# 0.0225f
C1169 xaa1.xa4.M0.D m2_4468_96284# 71.5f
C1170 xaa6.xg.XA1.MN0.D a_36172_53102# 0.00176f
C1171 a_36172_53454# a_37324_53454# 0.00133f
C1172 xaa1.xa4.M0.D m3_4788_74364# 0.0138f
C1173 li_4468_82684# li_4468_81884# 39.3f
C1174 xaa5.xb2_2.MN0.D a_29764_62158# 0.00263f
C1175 a_27244_62510# a_27244_62158# 0.0109f
C1176 xaa0.xa6.MN0.D xaa1.xa1.M0.D 8.17e-19
C1177 xaa1.xa2.M3.D PWRUP_1V8 0.00143f
C1178 AVDD a_5844_62366# 0.364f
C1179 xaa6.xd.XA7.MN1.G xaa6.xe.XA7.MN1.G 0.0108f
C1180 xaa6.xf.XA1.MN0.G a_36172_57326# 0.00148f
C1181 xaa6.xd.XA7.MP1.G xaa6.xe.XA7.MP1.G 0.00435f
C1182 xaa0.xa5.MN2.G xaa0.xa5.MN2.D 0.011f
C1183 a_36172_57678# xaa6.xg.XA7.MP1.G 2.36e-20
C1184 a_37324_57678# xaa6.xg.XA7.MN1.G 6.07e-19
C1185 PWRUP_1V8 a_34804_56270# 0.0079f
C1186 a_29764_57678# a_29764_57326# 0.0109f
C1187 xaa6.xg.XA7.MN1.D a_34804_57326# 1.31e-19
C1188 AVDD a_37324_56270# 0.362f
C1189 xaa6.xd.XA1.MN0.G xaa6.xe.XA1.MN0.D 0.00168f
C1190 a_2948_70022# li_4468_69404# 7.62e-20
C1191 xaa1.xa4.M0.D m1_4468_110684# 67.7f
C1192 xaa6.xg.XA7.MN1.D a_37324_53806# 0.0016f
C1193 a_31132_55918# xaa6.xe.XA5.MN0.G 0.0731f
C1194 a_244_53454# a_244_53102# 0.0109f
C1195 xaa1.xa4.M0.D m3_37668_90844# 0.074f
C1196 xaa3.xa7.MN0.D a_4692_62718# 0.00331f
C1197 xaa5.xa3.xb1_0.G a_28612_63566# 0.00581f
C1198 xaa4.xa2.M0.G xaa5.xa3.xb2_0.G 0.416f
C1199 a_28612_63918# a_29764_63918# 0.00133f
C1200 a_5844_63422# a_5844_63070# 0.0109f
C1201 xaa5.xb1.MN1.G a_29764_63566# 0.00513f
C1202 IBPSR_1U xaa1.xa2.M7.D 0.026f
C1203 m1_4468_114524# m2_4468_114524# 12.9f
C1204 a_26092_58030# a_27244_58030# 0.00133f
C1205 AVDD a_34804_57326# 0.00151f
C1206 m2_4468_96284# m3_37748_96604# 0.0138f
C1207 a_32284_56622# xaa6.xe.XA6.MN0.G 5.6e-19
C1208 xaa6.xf.XA1.MN0.G a_34804_55214# 0.00204f
C1209 xaa6.xd.XA7.MN1.G xaa6.xd.XA4.MP0.D 0.00941f
C1210 xaa6.xd.XA7.MP1.G xaa6.xd.XA4.MN0.D 0.056f
C1211 xaa6.xc.XA1.MN0.G a_28612_54862# 0.00209f
C1212 xaa1.xa4.M0.D li_4468_94204# 23f
C1213 PWRUP_1V8 a_34804_53806# 0.0737f
C1214 AVDD a_37324_53806# 0.405f
C1215 a_36172_54862# xaa6.xg.XA3.MN1.G 0.0723f
C1216 xaa6.xd.XA3.MP0.D xaa6.xd.XA3.MN0.D 0.00918f
C1217 CK_REF a_n908_52750# 4.33e-19
C1218 xaa1.xa4.M0.D m3_37748_108124# 0.111f
C1219 a_5844_57790# li_6204_57236# 5.99e-19
C1220 a_4692_57790# li_4836_56708# 9.91e-20
C1221 xaa3.xa1capd.B li_4980_56708# 0.0249f
C1222 xaa4.xa2.M0.G m3_13044_60468# 0.106f
C1223 li_4468_116444# li_4468_116284# 7.91f
C1224 a_356_70022# a_1220_70022# 0.071f
C1225 CK a_36172_58030# 4.94e-19
C1226 AVDD a_5844_60078# 0.364f
C1227 m2_4468_109724# m3_37668_110044# 0.0138f
C1228 xaa3.xa1capd.B a_5844_55150# 2.62e-19
C1229 xaa6.xg.XA7.MN1.D a_36172_56270# 0.012f
C1230 xaa6.xe.XA7.MN2.D a_31132_56974# 0.0494f
C1231 xaa3.xa1b.MN0.D a_4308_53678# 3.62e-19
C1232 IBPSR_1U xaa4.xa1.M4.D 0.026f
C1233 PWRUP_1V8 a_31132_55214# 0.00579f
C1234 xaa6.xe.XA7.MN1.D xaa6.xe.XA6.MN0.G 0.224f
C1235 xaa6.xf.XA1.MN0.G a_37324_56270# 1.11e-19
C1236 xaa6.xd.XA7.MP1.G xaa6.xd.XA6.MN0.D 0.056f
C1237 xaa6.xd.XA7.MN1.G xaa6.xd.XA6.MP0.D 0.0285f
C1238 xaa6.xc.XA7.MN1.D a_26092_55918# 0.00829f
C1239 AVDD a_33652_55214# 0.364f
C1240 a_33652_55566# a_33652_55214# 0.0109f
C1241 xaa1.xa4.M0.D m2_4468_97244# 71.5f
C1242 a_28612_53454# a_28612_53102# 0.0109f
C1243 xaa1.xa4.M0.D m3_4628_74364# 0.0276f
C1244 li_4468_106844# m1_4468_106844# 23f
C1245 xaa5.xb2_2.MN0.D a_28612_62158# 0.00224f
C1246 xaa3.xa1b.MN0.D a_4692_60782# 0.00455f
C1247 a_29764_62510# xaa5.xb2_1.MN0.D 0.0682f
C1248 xaa5.xa4.MN0.D xaa5.xa3.xb1_0.D 0.0638f
C1249 AVDD a_4692_62366# 0.00171f
C1250 m1_4468_80924# m2_4468_80924# 12.9f
C1251 xaa6.xf.XA7.MN1.D a_36172_57326# 1.31e-19
C1252 xaa6.xf.XA1.MN0.G a_34804_57326# 0.00134f
C1253 xaa0.xa5.MN2.G xaa0.xa5.MN0.D 0.22f
C1254 a_36172_57678# xaa6.xg.XA7.MN1.G 0.0736f
C1255 xaa6.xd.XA7.MN1.G xaa6.xd.XA7.MN0.D 0.0449f
C1256 AVDD a_36172_56270# 0.00151f
C1257 m2_4468_82844# m3_37748_83164# 0.0138f
C1258 xaa6.xd.XA1.MN0.G xaa6.xd.XA1.MN0.D 0.0147f
C1259 a_2948_70022# li_4468_70204# 6.88e-20
C1260 xaa1.xa4.M0.D m1_4468_111644# 67.7f
C1261 xaa6.xg.XA7.MN1.D a_36172_53806# 3.97e-20
C1262 xaa6.xf.XA7.MN1.G a_34804_54158# 0.0786f
C1263 xaa6.xf.XA1.MN0.G a_37324_53806# 1.11e-19
C1264 xaa6.xd.XA6.MN0.G a_29764_55566# 0.00224f
C1265 a_28612_54158# a_28612_53806# 0.0109f
C1266 xaa1.xa4.M0.D m3_4788_91644# 0.0138f
C1267 li_4468_99964# li_4468_99164# 39.3f
C1268 xaa5.xb3.MP1.D xaa5.xb2_3.MN0.D 7.69e-20
C1269 a_n908_63270# xaa1.xa2.M7.D 0.00155f
C1270 xaa5.xa3.xb1_0.G xaa5.xa3.xb2_0.G 1.05f
C1271 xaa5.xb1.MN1.G a_28612_63566# 9.6e-19
C1272 xaa4.xa2.M0.G a_29764_63918# 3.48e-19
C1273 PWRUP_1V8 a_31132_57326# 0.00561f
C1274 AVDD a_33652_57326# 0.364f
C1275 m2_4468_96284# m3_37668_96604# 0.0138f
C1276 xaa6.xd.XA7.MP1.G xaa6.xd.XA4.MP0.D 0.0615f
C1277 xaa6.xf.XA1.MN0.G a_33652_55214# 1.17e-19
C1278 a_36172_56622# a_36172_56270# 0.0109f
C1279 xaa6.xf.XA7.MN1.D a_34804_55214# 0.00558f
C1280 xaa6.xc.XA1.MN0.G a_27244_54862# 0.00257f
C1281 PWRUP_1V8 a_33652_53806# 0.0674f
C1282 AVDD a_36172_53806# 0.00156f
C1283 a_28612_54862# a_28612_54510# 0.0109f
C1284 xaa1.xa4.M0.D m3_37668_108124# 0.074f
C1285 a_5844_57790# li_6132_57236# 2e-19
C1286 xaa3.xa1capd.B li_4836_56708# 0.0139f
C1287 xaa4.xa2.M0.G m3_22620_61348# 0.0273f
C1288 xaa6.xg.XA5.MN0.G m1_37504_55818# 0.0386f
C1289 a_n940_70022# xaa1.xa3.D 0.0188f
C1290 CK a_34804_58030# 6.39e-19
C1291 AVDD a_4692_60078# 0.00171f
C1292 xaa3.xa1capd.B a_4692_55150# 1e-19
C1293 IBPSR_1U a_4308_53678# 0.0989f
C1294 PWRUP_1V8 a_29764_55214# 0.00579f
C1295 xaa6.xf.XA1.MN0.G a_36172_56270# 0.00193f
C1296 xaa4.xa4.M0.D xaa4.xa1.M8.D 0.218f
C1297 xaa6.xd.XA7.MP1.G xaa6.xd.XA6.MP0.D 0.0619f
C1298 xaa6.xd.XA1.MN0.G xaa6.xe.XA6.MN0.G 0.0171f
C1299 AVDD a_32284_55214# 0.364f
C1300 m2_4468_69404# m3_37748_69724# 0.0138f
C1301 xaa6.xe.XA5.MN0.G a_32284_54862# 0.0225f
C1302 xaa6.xe.XA6.MN0.G a_32284_54510# 0.00119f
C1303 xaa1.xa4.M0.D m2_4468_98204# 71.5f
C1304 xaa6.xf.XA1.MN0.D a_34804_53102# 0.00176f
C1305 a_34804_53454# a_36172_53454# 8.89e-19
C1306 xaa1.xa4.M0.D m3_37748_74524# 0.111f
C1307 li_4468_82844# li_4468_82684# 7.91f
C1308 a_26092_62510# a_26092_62158# 0.0109f
C1309 xaa0.xa6.MN0.D xaa1.xa1.M1.D 8.17e-19
C1310 a_28612_62510# xaa5.xb2_1.MN0.D 0.0674f
C1311 CK a_29764_62158# 3.97e-20
C1312 xaa1.xa2.M3.D xaa1.xa1.M8.D 0.00119f
C1313 xaa1.xa2.M4.D PWRUP_1V8 0.00107f
C1314 xaa6.xf.XA7.MN1.D a_34804_57326# 0.014f
C1315 xaa6.xd.XA7.MP1.G xaa6.xd.XA7.MN0.D 0.117f
C1316 a_28612_57678# a_28612_57326# 0.0109f
C1317 AVDD a_34804_56270# 0.00151f
C1318 m2_4468_82844# m3_37668_83164# 0.0138f
C1319 a_2948_70022# li_4468_70364# 3.68e-19
C1320 xaa1.xa4.M0.D m1_4468_112604# 67.7f
C1321 xaa6.xf.XA7.MP1.G a_34804_54158# 0.057f
C1322 xaa6.xf.XA7.MN1.G a_33652_54158# 0.0756f
C1323 a_29764_55918# xaa6.xd.XA5.MN0.G 0.0715f
C1324 xaa6.xf.XA1.MN0.G a_36172_53806# 0.00207f
C1325 xaa6.xd.XA6.MN0.G a_28612_55566# 0.0154f
C1326 xaa0.xa1.MP1.D a_244_53102# 0.00176f
C1327 a_n908_53454# a_n908_53102# 0.0109f
C1328 a_10092_54510# xaa4.xa1.M0.D 5.02e-20
C1329 xaa1.xa4.M0.D m3_4628_91644# 0.0276f
C1330 a_4692_63422# a_4692_63070# 0.0109f
C1331 xaa5.xa3.xb1_0.G a_29764_63918# 0.133f
C1332 xaa4.xa2.M0.G a_28612_63918# 0.0347f
C1333 xaa5.xb1.MN1.G xaa5.xa3.xb2_0.G 0.0625f
C1334 xaa3.xa7.MN0.D xaa3.xa6.MN0.D 0.128f
C1335 xaa0.xa6.MN0.D xaa1.xa2.M5.D 8.17e-19
C1336 m1_4468_115484# m2_4468_115484# 12.9f
C1337 PWRUP_1V8 a_29764_57326# 0.00567f
C1338 AVDD a_32284_57326# 0.364f
C1339 xaa6.xe.XA1.MN0.G a_34804_55214# 1.02e-19
C1340 xaa6.xf.XA7.MN1.D a_33652_55214# 0.00133f
C1341 xaa6.xc.XA7.MN1.D a_27244_54862# 0.00464f
C1342 xaa6.xc.XA6.MN0.D xaa6.xc.XA6.MP0.D 0.00918f
C1343 xaa6.xc.XA1.MN0.G a_26092_54862# 4.77e-19
C1344 xaa1.xa4.M0.D li_4468_95164# 23f
C1345 PWRUP_1V8 a_32284_53806# 0.0658f
C1346 AVDD a_34804_53806# 0.00156f
C1347 CK_REF a_n908_53102# 8.56e-19
C1348 a_34804_54862# xaa6.xf.XA3.MN0.D 0.00176f
C1349 xaa1.xa4.M0.D m3_4788_108924# 0.0138f
C1350 xaa3.xa1capd.B li_6204_57236# 0.118f
C1351 xaa6.xg.XA5.MN0.D m1_37504_55818# 0.0453f
C1352 xaa4.xa2.M0.G m3_22548_61348# 0.0137f
C1353 li_4468_117244# li_4468_116444# 39.3f
C1354 a_2948_74698# xaa1.xa3.D 1.91e-21
C1355 xaa1.xa4.M0.D a_2948_70022# 0.00777f
C1356 li_4468_84764# m1_4468_84764# 23f
C1357 PWRUP_1V8 xaa1.xa1.M0.D 4.28e-19
C1358 xaa1.xa1.M8.D xaa1.xb1.M0.D 0.099f
C1359 CK a_33652_58030# 2.89e-19
C1360 xaa0.xa2a.MN0.D xaa1.xa1.M3.D 0.00394f
C1361 AVDD xaa1.xb1.M0.D 0.085f
C1362 xaa3.xa1capd.B a_5844_55502# 7.03e-19
C1363 IBPSR_1U a_244_52750# 0.00162f
C1364 xaa6.xf.XA1.MN0.G a_34804_56270# 0.00204f
C1365 CK xaa6.xg.XA3.MN1.G 0.0676f
C1366 xaa6.xd.XA1.MN0.G xaa6.xd.XA6.MN0.G 0.0112f
C1367 xaa6.xd.XA7.MN2.D a_29764_56974# 0.0494f
C1368 AVDD a_31132_55214# 0.00151f
C1369 m2_4468_69404# m3_37668_69724# 0.0138f
C1370 xaa6.xg.XA7.MN1.G a_37324_52750# 0.00141f
C1371 xaa6.xe.XA5.MN0.G a_31132_54862# 0.033f
C1372 a_32284_55566# a_32284_55214# 0.0109f
C1373 xaa1.xa4.M0.D m2_4468_99164# 71.5f
C1374 a_4308_53678# xbb1.xa3.M0.D 5.02e-20
C1375 a_27244_53454# a_27244_53102# 0.0109f
C1376 xaa4.xa1.M2.D a_10092_52750# 2.99e-19
C1377 a_37324_56974# m1_37504_55818# 2.34e-19
C1378 xaa1.xa4.M0.D m3_37668_74524# 0.074f
C1379 xaa5.xa3.xb2_0.G a_26092_61102# 0.00183f
C1380 IBPSR_1U xaa1.xa1.M3.D 0.026f
C1381 xaa4.xa2.M0.G a_29764_61102# 2.68e-19
C1382 xaa5.xa3.xb2_0.D a_27244_62158# 0.0318f
C1383 AVDD xaa3.xa5a.MN0.D 1.12f
C1384 m1_4468_81884# m2_4468_81884# 12.9f
C1385 a_34804_57678# xaa6.xf.XA7.MN0.D 0.00176f
C1386 xaa6.xf.XA7.MN1.D a_33652_57326# 0.00337f
C1387 xaa6.xe.XA1.MN0.G a_34804_57326# 0.0662f
C1388 xaa0.xa5.MN2.G a_n908_56622# 0.00164f
C1389 PWRUP_1V8 a_31132_56270# 0.00783f
C1390 xaa6.xd.XA7.MP1.G xaa6.xd.XA7.MN1.G 0.537f
C1391 AVDD a_33652_56270# 0.363f
C1392 xaa6.xc.XA1.MN0.G xaa6.xd.XA1.MN0.D 2.73e-19
C1393 a_2948_70022# li_4468_71164# 1.04e-19
C1394 xaa1.xa3.D li_4468_70204# 0.00464f
C1395 xaa1.xa4.M0.D m1_4468_113564# 67.7f
C1396 xaa6.xf.XA7.MP1.G a_33652_54158# 0.0545f
C1397 xaa6.xf.XA7.MN1.G a_32284_54158# 7.1e-20
C1398 a_28612_55918# xaa6.xd.XA5.MN0.G 0.0674f
C1399 xaa6.xf.XA1.MN0.G a_34804_53806# 0.0032f
C1400 xaa6.xg.XA6.MN0.G xaa6.xg.XA5.MN0.G 0.0629f
C1401 a_n908_53454# a_244_53454# 0.00133f
C1402 a_27244_54158# a_27244_53806# 0.0109f
C1403 xaa1.xa4.M0.D m3_37748_91804# 0.111f
C1404 li_4468_100124# li_4468_99964# 7.91f
C1405 xaa3.xa8.MP0.D a_5844_63070# 0.00176f
C1406 xaa5.xb3.MP1.D a_28612_63214# 1.02e-19
C1407 xaa5.xa3.xb1_0.G a_28612_63918# 0.0958f
C1408 xaa5.xb1.MN1.G a_29764_63918# 0.00811f
C1409 xaa4.xa4.M0.D xaa0.xa5.MN2.G 5.35e-20
C1410 AVDD a_31132_57326# 0.00151f
C1411 a_34804_56622# a_34804_56270# 0.0109f
C1412 xaa6.xe.XA1.MN0.G a_33652_55214# 0.00196f
C1413 xaa6.xc.XA7.MN1.D a_26092_54862# 0.00652f
C1414 PWRUP_1V8 a_31132_53806# 0.0753f
C1415 AVDD a_33652_53806# 0.406f
C1416 xaa1.xa4.M0.D m3_4628_108924# 0.0276f
C1417 xaa0.xa1.MN0.D a_244_52750# 5.1e-20
C1418 a_27244_54862# a_27244_54510# 0.0109f
C1419 CK_REF a_244_53454# 0.0674f
C1420 xaa3.xa1capd.B li_6132_57236# 0.0319f
C1421 xaa4.xa2.M0.G m3_13116_61524# 0.0634f
C1422 a_28612_61102# a_29764_61102# 0.00133f
C1423 CK a_32284_58030# 9.38e-19
C1424 xaa0.xa2a.MN0.D a_640_60806# 0.0705f
C1425 AVDD xaa3.xa3a.MN0.D 1.12f
C1426 IBPSR_1U a_n908_52750# 0.00131f
C1427 xaa6.xf.XA7.MN1.D a_34804_56270# 0.012f
C1428 xaa6.xf.XA1.MN0.G a_33652_56270# 1.17e-19
C1429 xaa6.xd.XA7.MN1.D xaa6.xd.XA6.MN0.G 0.224f
C1430 xaa3.xa1capd.B a_4692_55502# 2.12e-19
C1431 xaa6.xg.XA7.MN0.G xaa6.xg.XA7.MN2.D 0.00981f
C1432 AVDD a_29764_55214# 0.00151f
C1433 xaa1.xa4.M0.D m2_4468_100124# 71.5f
C1434 xaa1.xa4.M0.D m3_4788_75324# 0.0138f
C1435 a_4308_53678# xbb1.xa3.M1.D 6.46e-20
C1436 a_33652_53454# a_34804_53454# 0.00133f
C1437 a_37324_56974# m1_37504_57930# 0.00375f
C1438 li_4468_83644# li_4468_82844# 39.3f
C1439 li_4468_107804# m1_4468_107804# 23f
C1440 IBPSR_1U a_640_60806# 6.96e-19
C1441 xaa4.xa2.M0.G a_28612_61102# 0.0189f
C1442 xaa1.xa3.D a_640_59750# 5.02e-20
C1443 a_27244_62510# xaa5.xa3.xb1_0.D 0.0673f
C1444 xaa5.xa3.xb2_0.D a_26092_62158# 0.0571f
C1445 xaa1.xa2.M4.D xaa1.xa1.M8.D 8.35e-19
C1446 a_33652_57678# xaa6.xf.XA7.MN0.D 0.00176f
C1447 a_34804_57678# xaa6.xf.XA7.MN1.G 0.072f
C1448 xaa6.xe.XA1.MN0.G a_33652_57326# 0.0858f
C1449 xaa0.xa5.MN2.G xaa0.xa3.MN1.G 0.116f
C1450 PWRUP_1V8 a_29764_56270# 0.0079f
C1451 a_27244_57678# a_27244_57326# 0.0109f
C1452 AVDD a_32284_56270# 0.363f
C1453 xaa1.xa4.M0.D m1_4468_114524# 67.7f
C1454 a_2948_70022# li_4468_71324# 3.68e-19
C1455 xaa6.xc.XA1.MN0.G xaa6.xc.XA1.MN0.D 0.0357f
C1456 xaa6.xg.XA6.MN0.G xaa6.xg.XA5.MN0.D 0.00862f
C1457 xaa6.xf.XA7.MN1.D a_34804_53806# 3.97e-20
C1458 xaa6.xf.XA1.MN0.G a_33652_53806# 1.35e-19
C1459 xaa6.xc.XA6.MN0.G a_27244_55566# 0.0154f
C1460 a_37324_58030# m1_37504_57930# 0.00743f
C1461 xaa0.xa1.MP1.D a_244_53454# 0.0494f
C1462 xaa1.xa4.M0.D m3_37668_91804# 0.074f
C1463 xaa6.xg.XA3.MP0.D m1_37504_55818# 8.78e-20
C1464 xaa1.xa2.M8.D xaa1.xa2.M7.D 0.0488f
C1465 xaa5.xa3.xb1_0.G xaa4.xa2.M0.G 0.414f
C1466 xaa5.xb1.MN1.G a_28612_63918# 0.0032f
C1467 xaa3.xa7.MN0.D a_5844_63070# 0.022f
C1468 xaa0.xa6.MN0.D xaa1.xa2.M6.D 8.17e-19
C1469 m1_4468_116444# m2_4468_116444# 12.9f
C1470 a_4692_57790# a_5844_57790# 0.00133f
C1471 AVDD a_29764_57326# 0.00151f
C1472 a_28612_56622# xaa6.xd.XA6.MN0.G 5.6e-19
C1473 xaa6.xe.XA1.MN0.G a_32284_55214# 0.00207f
C1474 xaa1.xa4.M0.D li_4468_96124# 23f
C1475 PWRUP_1V8 a_29764_53806# 0.0737f
C1476 xaa6.xc.XA7.MP1.G xaa6.xc.XA4.MP0.D 0.0615f
C1477 AVDD a_32284_53806# 0.406f
C1478 xaa1.xa4.M0.D m3_37748_109084# 0.111f
C1479 xaa6.xc.XA3.MN0.D xaa6.xc.XA3.MP0.D 0.00918f
C1480 xaa0.xa1.MN0.D a_n908_52750# 1.28e-19
C1481 a_244_53806# a_244_53454# 0.0109f
C1482 a_33652_54862# xaa6.xf.XA3.MP0.D 0.00176f
C1483 CK_REF a_n908_53454# 0.0658f
C1484 xaa4.xa2.M0.G m3_13044_61524# 0.106f
C1485 li_4468_117404# li_4468_117244# 7.91f
C1486 xaa1.xa4.M0.D xaa1.xa3.D 4f
C1487 xaa0.xa2a.MN0.D xaa1.xa1.M4.D 0.00573f
C1488 xaa1.xa1.M8.D xaa1.xa1.M0.D 8.76e-19
C1489 PWRUP_1V8 xaa1.xa1.M1.D 5.67e-19
C1490 AVDD xaa1.xa1.M0.D 5.56e-19
C1491 m2_4468_110684# m3_37748_111004# 0.0138f
C1492 xaa6.xc.XA7.MP1.G xaa6.xc.XA6.MP0.D 0.0619f
C1493 IBPSR_1U a_244_53102# 4.86e-19
C1494 PWRUP_1V8 a_26092_55214# 0.00572f
C1495 xaa6.xf.XA7.MN1.D a_33652_56270# 0.00378f
C1496 xaa6.xe.XA1.MN0.G a_34804_56270# 1.02e-19
C1497 xaa6.xc.XA1.MN0.G xaa6.xd.XA6.MN0.G 0.0181f
C1498 AVDD a_28612_55214# 0.364f
C1499 xaa6.xd.XA5.MN0.G a_29764_54862# 0.033f
C1500 xaa4.xa2.M0.D a_10092_54510# 0.00733f
C1501 a_31132_55566# a_31132_55214# 0.0109f
C1502 xaa6.xg.XA5.MN0.G xaa6.xg.XA4.MN0.G 0.0564f
C1503 a_2948_70022# m1_4468_69404# 2.28e-19
C1504 xaa1.xa4.M0.D m2_4468_101084# 71.5f
C1505 xaa1.xa4.M0.D m3_4628_75324# 0.0276f
C1506 a_4308_53678# xbb1.xa3.M2.D 8.62e-20
C1507 a_26092_53454# a_26092_53102# 0.0109f
C1508 xaa5.xb1.MN1.G a_29764_61102# 0.0732f
C1509 IBPSR_1U xaa1.xa1.M4.D 0.026f
C1510 xaa4.xa2.M0.G a_27244_61102# 5.56e-19
C1511 xaa5.xb2_2.MN0.D xaa5.xb2_1.MN0.D 0.197f
C1512 a_26092_62510# xaa5.xa3.xb1_0.D 0.0728f
C1513 a_27244_62510# xaa5.xa4.MN0.D 0.0215f
C1514 a_28612_62510# a_29764_62510# 0.00133f
C1515 xaa1.xa2.M3.D a_n908_61510# 1.81e-19
C1516 CK a_26092_62158# 3.16e-19
C1517 xaa1.xa2.M5.D PWRUP_1V8 8.33e-19
C1518 AVDD a_5844_62718# 0.388f
C1519 m1_4468_82844# m2_4468_82844# 12.9f
C1520 a_33652_57678# xaa6.xf.XA7.MN1.G 5.46e-19
C1521 a_34804_57678# xaa6.xf.XA7.MP1.G 2.36e-20
C1522 xaa6.xe.XA1.MN0.G a_32284_57326# 0.00236f
C1523 xaa6.xc.XA7.MP1.G xaa6.xd.XA7.MN1.G 1.74e-19
C1524 AVDD a_31132_56270# 0.00151f
C1525 xaa1.xa4.M0.D m1_4468_115484# 67.7f
C1526 xaa1.xa3.D li_4468_71164# 0.00464f
C1527 a_2948_70022# li_4468_72124# 1.04e-19
C1528 a_36172_55918# a_37324_55918# 0.00133f
C1529 a_27244_55918# xaa6.xc.XA5.MN0.G 0.0658f
C1530 xaa6.xf.XA7.MN1.D a_33652_53806# 0.0016f
C1531 xaa6.xe.XA1.MN0.G a_34804_53806# 1.11e-19
C1532 xaa6.xc.XA6.MN0.G a_26092_55566# 0.00224f
C1533 a_26092_54158# a_26092_53806# 0.0109f
C1534 xaa1.xa4.M0.D m3_4788_92604# 0.0138f
C1535 li_4468_100924# li_4468_100124# 39.3f
C1536 xaa1.xa4.M0.G xaa3.xa5a.MN0.D 5.72e-20
C1537 xaa5.xb1.MN1.G xaa4.xa2.M0.G 0.132f
C1538 xaa3.xa7.MN0.D a_4692_63070# 0.057f
C1539 PWRUP_1V8 a_26092_57326# 0.00579f
C1540 xaa3.xa1capd.B a_5844_57790# 0.0766f
C1541 AVDD a_28612_57326# 0.364f
C1542 m2_4468_97244# m3_37748_97564# 0.0138f
C1543 xaa6.xe.XA1.MN0.G a_31132_55214# 1.06e-19
C1544 a_33652_56622# a_33652_56270# 0.0109f
C1545 xaa6.xe.XA7.MN1.D a_32284_55214# 0.00133f
C1546 PWRUP_1V8 a_28612_53806# 0.0674f
C1547 xaa6.xc.XA7.MP1.G xaa6.xc.XA4.MN0.D 0.056f
C1548 xaa6.xc.XA7.MN1.G xaa6.xc.XA4.MP0.D 0.00941f
C1549 AVDD a_31132_53806# 0.00156f
C1550 xaa1.xa4.M0.D m3_37668_109084# 0.074f
C1551 CK_REF xaa0.xa1.MP1.D 0.00999f
C1552 xaa0.xa1.MN0.D a_244_53102# 1.28e-19
C1553 a_26092_54862# a_26092_54510# 0.0109f
C1554 a_2084_74698# xaa1.xa3.D 0.00296f
C1555 li_4468_85724# m1_4468_85724# 23f
C1556 xaa0.xa2a.MN0.D xaa1.xb2.M7.D 0.0157f
C1557 xaa1.xa1.M5.D xaa1.xa1.M4.D 0.0488f
C1558 xaa1.xa1.M8.D a_640_60278# 0.182f
C1559 a_27244_61102# a_28612_61102# 8.89e-19
C1560 AVDD a_640_60278# 0.385f
C1561 m2_4468_110684# m3_37668_111004# 0.0138f
C1562 IBPSR_1U a_n908_53102# 4.86e-19
C1563 xaa6.xc.XA7.MN1.G xaa6.xc.XA6.MP0.D 0.0285f
C1564 xaa6.xc.XA7.MP1.G xaa6.xc.XA6.MN0.D 0.056f
C1565 xaa6.xe.XA1.MN0.G a_33652_56270# 0.00211f
C1566 xaa6.xc.XA1.MN0.G xaa6.xc.XA6.MN0.G 0.0125f
C1567 AVDD a_27244_55214# 0.364f
C1568 xaa6.xd.XA5.MN0.G a_28612_54862# 0.0225f
C1569 xaa6.xd.XA6.MN0.G a_28612_54510# 0.00119f
C1570 xaa6.xg.XA5.MN0.G a_37324_55214# 0.00301f
C1571 a_244_53806# CK_REF 0.0658f
C1572 a_37324_55566# xaa6.xg.XA4.MP0.D 0.00176f
C1573 a_2948_70022# m1_4468_70204# 1.79e-19
C1574 xaa1.xa4.M0.D m2_4468_102044# 71.5f
C1575 xaa1.xa4.M0.D m3_37748_75484# 0.111f
C1576 a_32284_53454# a_33652_53454# 8.89e-19
C1577 xaa6.xe.XA1.MN0.D a_31132_53102# 0.00176f
C1578 li_4468_83804# li_4468_83644# 7.91f
C1579 xaa0.xa6.MN0.D xaa1.xa1.M2.D 8.17e-19
C1580 xaa1.xa3.D xaa4.xa4.M0.D 0.0439f
C1581 xaa5.xb1.MN1.G a_28612_61102# 0.0658f
C1582 xaa5.xa3.xb1_0.G a_27244_61102# 2.6e-19
C1583 AVDD a_4692_62718# 0.00171f
C1584 a_26092_62510# xaa5.xa4.MN0.D 0.0215f
C1585 xaa6.xe.XA1.MN0.G a_31132_57326# 1.06e-19
C1586 a_33652_57678# xaa6.xf.XA7.MP1.G 0.071f
C1587 xaa6.xe.XA7.MN1.D a_32284_57326# 0.00337f
C1588 xaa0.xa5.MN2.G a_n908_56974# 4.46e-19
C1589 xaa6.xc.XA7.MN1.G xaa6.xd.XA7.MN1.G 0.31f
C1590 xaa6.xc.XA7.MP1.G xaa6.xd.XA7.MP1.G 0.00435f
C1591 xaa6.xd.XA1.MN0.G a_33652_57326# 2.93e-19
C1592 a_26092_57678# a_26092_57326# 0.0109f
C1593 AVDD a_29764_56270# 0.00151f
C1594 m2_4468_83804# m3_37748_84124# 0.0138f
C1595 xaa1.xa4.M0.D m1_4468_116444# 67.7f
C1596 a_2948_70022# li_4468_72284# 2e-19
C1597 xaa6.xe.XA7.MP1.G a_32284_54158# 0.0545f
C1598 xaa6.xe.XA7.MN1.G a_33652_54158# 7.1e-20
C1599 xaa6.xf.XA6.MN0.G xaa6.xf.XA5.MN0.G 0.27f
C1600 a_26092_55918# xaa6.xc.XA5.MN0.G 0.0731f
C1601 xaa6.xe.XA1.MN0.G a_33652_53806# 0.00209f
C1602 xaa6.xg.XA3.MN1.G xaa6.xg.XA1.MN0.D 0.122f
C1603 xaa1.xa4.M0.D m3_4628_92604# 0.0276f
C1604 a_4692_63774# xaa3.xa6.MN0.D 1.73e-19
C1605 xaa5.xb1.MN1.G xaa5.xa3.xb1_0.G 0.194f
C1606 m1_4468_117404# m2_4468_117404# 12.9f
C1607 PWRUP_1V8 xaa6.xg.XA7.MN0.D 0.0493f
C1608 a_5844_58142# a_5844_57790# 0.0109f
C1609 xaa3.xa1capd.B a_4692_57790# 0.0913f
C1610 AVDD a_27244_57326# 0.364f
C1611 m2_4468_97244# m3_37668_97564# 0.0138f
C1612 xaa6.xg.XA7.MP1.G a_37324_55566# 0.0292f
C1613 a_27244_56622# xaa6.xc.XA6.MN0.G 5.6e-19
C1614 xaa6.xe.XA7.MN1.D a_31132_55214# 0.00558f
C1615 a_4692_55854# a_5844_55854# 0.00133f
C1616 xaa0.xa2a.MN0.D a_244_53454# 5.27e-19
C1617 xaa6.xd.XA1.MN0.G a_32284_55214# 1.11e-19
C1618 xaa1.xa4.M0.D li_4468_97084# 23f
C1619 PWRUP_1V8 a_27244_53806# 0.0658f
C1620 xaa6.xc.XA7.MN1.G xaa6.xc.XA4.MN0.D 1.09e-19
C1621 AVDD a_29764_53806# 0.00156f
C1622 xaa1.xa4.M0.D m3_4788_109884# 0.0138f
C1623 a_n908_53806# a_n908_53454# 0.0109f
C1624 a_244_53806# xaa0.xa1.MP1.D 0.00176f
C1625 a_32284_54862# xaa6.xe.XA3.MP0.D 0.00176f
C1626 xaa0.xa1.MN0.D a_n908_53102# 0.00385f
C1627 li_4468_118204# li_4468_117404# 39.3f
C1628 a_n76_72222# a_788_72222# 0.107f
C1629 xaa1.xa1.M8.D xaa1.xa1.M1.D 0.00115f
C1630 xaa6.xe.XA1.MN0.G a_32284_56270# 0.00207f
C1631 xaa6.xc.XA7.MN1.D xaa6.xc.XA6.MN0.G 0.224f
C1632 xaa6.xc.XA7.MN1.G xaa6.xc.XA6.MN0.D 0.0158f
C1633 xaa6.xc.XA7.MN2.D a_26092_56974# 0.0494f
C1634 AVDD a_26092_55214# 0.00159f
C1635 m2_4468_70364# m3_37748_70684# 0.0138f
C1636 xaa6.xg.XA5.MN0.G a_36172_55214# 0.0155f
C1637 a_n908_53806# CK_REF 0.0725f
C1638 a_29764_55566# a_29764_55214# 0.0109f
C1639 a_2948_70022# m1_4468_70364# 0.00161f
C1640 xaa1.xa4.M0.D m2_4468_103004# 71.5f
C1641 xaa6.xf.XA7.MN1.G a_34804_52750# 2.64e-19
C1642 xaa1.xa4.M0.D m3_37668_75484# 0.074f
C1643 xbb1.xa3.M5.D xbb1.xa3.M4.D 0.0488f
C1644 li_4468_108764# m1_4468_108764# 23f
C1645 xaa5.xa3.xb1_0.G a_26092_61102# 0.173f
C1646 xaa5.xa3.xb2_0.D xaa5.xa3.xb1_0.D 0.607f
C1647 CK xaa5.xb2_1.MN0.D 7.29e-20
C1648 a_27244_62510# a_28612_62510# 8.89e-19
C1649 xaa1.xa2.M4.D a_n908_61510# 1.21e-19
C1650 xaa1.xa2.M5.D xaa1.xa1.M8.D 6.17e-19
C1651 xaa1.xa2.M6.D PWRUP_1V8 6.63e-19
C1652 m1_4468_83804# m2_4468_83804# 12.9f
C1653 xaa6.xe.XA7.MN1.D a_31132_57326# 0.014f
C1654 xaa6.xc.XA7.MN1.G xaa6.xd.XA7.MP1.G 1.74e-19
C1655 xaa6.xd.XA1.MN0.G a_32284_57326# 0.081f
C1656 xaa6.xc.XA7.MP1.G xaa6.xc.XA7.MN0.D 0.117f
C1657 PWRUP_1V8 a_26092_56270# 0.00776f
C1658 AVDD a_28612_56270# 0.363f
C1659 m2_4468_83804# m3_37668_84124# 0.0138f
C1660 xaa1.xa4.M0.D m1_4468_117404# 67.7f
C1661 xaa1.xa3.D li_4468_72124# 0.00464f
C1662 a_2948_70022# li_4468_73084# 1.76e-20
C1663 a_34804_55918# a_36172_55918# 8.89e-19
C1664 xaa6.xe.XA7.MP1.G a_31132_54158# 0.057f
C1665 xaa6.xe.XA7.MN1.G a_32284_54158# 0.074f
C1666 xaa6.xe.XA1.MN0.G a_32284_53806# 0.0044f
C1667 xaa1.xa4.M0.D m3_37748_92764# 0.111f
C1668 li_4468_101084# li_4468_100924# 7.91f
C1669 xaa3.xa9.MN0.D xaa3.xa6.MN0.D 5.43e-20
C1670 IBPSR_1U xaa4.xa2.M0.G 0.0369f
C1671 xaa0.xa6.MN0.D xaa1.xa2.M7.D 8.17e-19
C1672 PWRUP_1V8 xaa6.xg.XA7.MP1.G 0.124f
C1673 AVDD a_26092_57326# 0.00159f
C1674 xaa3.xa1b.MN0.D a_5844_55854# 0.0901f
C1675 xaa6.xg.XA7.MP1.G a_36172_55566# 0.098f
C1676 xaa6.xg.XA7.MN1.G a_37324_55566# 0.00742f
C1677 a_32284_56622# a_32284_56270# 0.0109f
C1678 CK a_37324_53454# 0.0662f
C1679 xaa0.xa2a.MN0.D a_n908_53454# 8.92e-20
C1680 xaa6.xd.XA1.MN0.G a_31132_55214# 0.00193f
C1681 a_36172_57326# xaa6.xg.XA5.MN0.G 6.98e-20
C1682 PWRUP_1V8 a_26092_53806# 0.0752f
C1683 a_5844_56206# a_5844_55854# 0.0109f
C1684 AVDD a_28612_53806# 0.406f
C1685 xaa1.xa4.M0.D m3_4628_109884# 0.0276f
C1686 xaa0.xa1.MN2.D a_n908_53454# 0.00176f
C1687 xaa0.xa1.MN0.D a_244_53454# 0.00328f
C1688 xaa3.xa2.MN0.D li_4980_58996# 7.61e-20
C1689 a_26092_61102# a_27244_61102# 0.00133f
C1690 a_640_61158# a_640_60806# 0.0109f
C1691 a_n908_61510# xaa1.xa1.M0.D 5.02e-20
C1692 xaa4.xa2.M0.G a_11712_57502# 0.0188f
C1693 AVDD a_5844_60430# 0.388f
C1694 xaa6.xe.XA1.MN0.G a_31132_56270# 1.06e-19
C1695 PWRUP_1V8 xaa6.xg.XA4.MN0.D 0.00353f
C1696 xaa6.xe.XA7.MN1.D a_32284_56270# 0.00378f
C1697 xaa0.xa5.MN2.G xaa6.xc.XA6.MN0.G 0.00663f
C1698 xaa6.xg.XA7.MN0.D a_37324_56622# 0.0217f
C1699 a_37324_57326# a_37324_56974# 0.0109f
C1700 xaa0.xa2a.MN0.D CK_REF 0.00151f
C1701 AVDD a_10092_55038# 0.0011f
C1702 m2_4468_70364# m3_37668_70684# 0.0138f
C1703 xaa6.xc.XA5.MN0.G a_27244_54862# 0.0225f
C1704 xaa6.xc.XA6.MN0.G a_27244_54510# 0.00119f
C1705 a_n908_53806# a_244_53806# 0.00133f
C1706 a_37324_55566# xaa6.xg.XA4.MP1.G 0.0658f
C1707 a_36172_55566# xaa6.xg.XA4.MN0.D 0.00176f
C1708 xaa0.xa1.MN2.D CK_REF 0.0111f
C1709 a_2948_70022# m1_4468_71164# 1.79e-19
C1710 xaa1.xa3.D m1_4468_70204# 12.9f
C1711 xaa1.xa4.M0.D m2_4468_103964# 71.5f
C1712 xaa6.xf.XA7.MN1.G a_33652_52750# 0.00154f
C1713 xaa1.xa4.M0.D m3_4788_76284# 0.0138f
C1714 a_31132_53454# a_32284_53454# 0.00133f
C1715 xaa6.xd.XA1.MN0.D a_29764_53102# 0.00176f
C1716 li_4468_84604# li_4468_83804# 39.3f
C1717 xaa5.xa3.xb2_0.D xaa5.xa4.MN0.D 0.0773f
C1718 CK xaa5.xa3.xb1_0.D 0.00109f
C1719 xaa5.xb2_2.MN0.D a_29764_62510# 0.126f
C1720 AVDD xaa3.xa6.MN0.D 0.724f
C1721 xaa6.xc.XA7.MN1.G xaa6.xc.XA7.MN0.D 0.0449f
C1722 xaa6.xd.XA1.MN0.G a_31132_57326# 0.0689f
C1723 AVDD a_27244_56270# 0.363f
C1724 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MN0.D 0.336f
C1725 a_32284_57678# xaa6.xe.XA7.MN0.D 0.00176f
C1726 xaa6.xe.XA7.MN1.D a_29764_57326# 1.31e-19
C1727 xaa6.xe.XA6.MN0.G xaa6.xe.XA5.MN0.G 0.27f
C1728 xaa6.xe.XA7.MN1.G a_31132_54158# 0.0802f
C1729 xaa6.xe.XA7.MN1.D a_32284_53806# 0.0016f
C1730 xaa6.xe.XA1.MN0.G a_31132_53806# 0.00318f
C1731 xaa1.xa4.M0.D m3_37668_92764# 0.074f
C1732 xaa1.xa4.M0.G a_4692_62718# 5.18e-20
C1733 a_4692_58142# a_4692_57790# 0.0109f
C1734 a_5844_58142# xaa3.xa1capd.B 0.0658f
C1735 xaa3.xa2.MN0.D a_5844_57790# 0.00224f
C1736 a_26092_60750# xaa0.xa5.MN2.G 3.82e-19
C1737 PWRUP_1V8 xaa6.xg.XA7.MN1.G 0.275f
C1738 xaa3.xa1b.MN0.D a_4692_55854# 0.124f
C1739 AVDD xaa6.xg.XA7.MN0.D 0.485f
C1740 xaa6.xg.XA7.MN1.G a_36172_55566# 3.45e-19
C1741 a_33652_56974# xaa6.xf.XA6.MN0.G 2.34e-19
C1742 CK a_36172_53454# 0.0717f
C1743 xaa0.xa2a.MN0.D xaa0.xa1.MP1.D 9.65e-20
C1744 xaa6.xd.XA1.MN0.G a_29764_55214# 0.00204f
C1745 xaa1.xa4.M0.D li_4468_98044# 23f
C1746 xaa6.xg.XA7.MN1.D xaa6.xg.XA4.MP0.D 0.00426f
C1747 AVDD a_27244_53806# 0.406f
C1748 xaa1.xa4.M0.D m3_37748_110044# 0.111f
C1749 a_31132_54862# xaa6.xe.XA3.MN0.D 0.00176f
C1750 xaa0.xa1.MN0.D a_n908_53454# 0.0799f
C1751 xaa3.xa2.MN0.D li_4836_58996# 4.62e-19
C1752 xaa1.xa4.M0.D a_1652_72222# 2.87e-19
C1753 a_n508_70022# a_356_70022# 0.071f
C1754 li_4468_86684# m1_4468_86684# 23f
C1755 xaa5.xb1.MN0.D a_29764_61102# 0.0492f
C1756 PWRUP_1V8 xaa1.xa1.M2.D 5.67e-19
C1757 AVDD a_4692_60430# 0.00171f
C1758 xaa6.xe.XA7.MN1.D a_31132_56270# 0.012f
C1759 IBPSR_1U xaa0.xa1.MP1.D 1.76e-20
C1760 xaa6.xg.XA7.MP1.G a_37324_56622# 0.029f
C1761 xaa6.xd.XA1.MN0.G a_32284_56270# 2.6e-19
C1762 xaa4.xa4.M0.D a_10092_55566# 0.00541f
C1763 xaa6.xg.XA7.MN0.D a_36172_56622# 1.28e-19
C1764 xaa0.xa2a.MN0.D a_244_53806# 8.96e-19
C1765 AVDD xaa6.xg.XA4.MP0.D 0.159f
C1766 xaa0.xa1.MN2.S a_n908_53454# 0.0293f
C1767 xaa6.xc.XA5.MN0.G a_26092_54862# 0.033f
C1768 xaa0.xa1.MN0.D CK_REF 0.202f
C1769 a_28612_55566# a_28612_55214# 0.0109f
C1770 a_2948_70022# m1_4468_71324# 0.00161f
C1771 xaa1.xa4.M0.D m2_4468_104924# 71.5f
C1772 xaa1.xa4.M0.D m3_4628_76284# 0.0276f
C1773 xaa4.xa1.M1.D xaa4.xa1.M0.D 0.0488f
C1774 xaa4.xa2.M0.G xaa5.xb1.MN0.D 1.92e-19
C1775 CK xaa5.xa4.MN0.D 0.0476f
C1776 xaa5.xb2_2.MN0.D a_28612_62510# 0.0878f
C1777 a_26092_62510# a_27244_62510# 0.00133f
C1778 xaa1.xa2.M6.D xaa1.xa1.M8.D 4.74e-19
C1779 m1_4468_84764# m2_4468_84764# 12.9f
C1780 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MP1.G 0.314f
C1781 xaa6.xd.XA7.MN1.D a_31132_57326# 1.31e-19
C1782 xaa6.xd.XA1.MN0.G a_29764_57326# 0.00134f
C1783 AVDD a_26092_56270# 0.00159f
C1784 PWRUP_1V8 xaa6.xg.XA6.MN0.D 0.00353f
C1785 a_32284_57678# xaa6.xe.XA7.MP1.G 0.0694f
C1786 xaa6.xc.XA7.MN1.G xaa6.xc.XA7.MP1.G 0.537f
C1787 a_31132_57678# xaa6.xe.XA7.MN0.D 0.00176f
C1788 a_33652_55918# a_34804_55918# 0.00133f
C1789 a_37324_56270# xaa6.xg.XA5.MN0.D 2.54e-19
C1790 xaa6.xe.XA7.MN1.D a_31132_53806# 3.97e-20
C1791 xaa0.xa1.MN2.S CK_REF 0.104f
C1792 a_36172_56270# xaa6.xg.XA5.MN0.G 0.00131f
C1793 xaa6.xd.XA1.MN0.G a_32284_53806# 1.11e-19
C1794 a_36172_54158# a_37324_54158# 0.00133f
C1795 xaa4.xa1.M5.D xaa4.xa1.M4.D 0.0488f
C1796 xaa1.xa4.M0.D m3_4788_93564# 0.0138f
C1797 li_4468_101884# li_4468_101084# 39.3f
C1798 a_4692_64126# xaa3.xa6.MN0.D 1.76e-20
C1799 a_4692_58142# xaa3.xa1capd.B 0.0728f
C1800 xaa3.xa2.MN0.D a_4692_57790# 0.00346f
C1801 PWRUP_1V8 xaa6.xf.XA7.MN0.D 0.0493f
C1802 IBPSR_1U a_4692_55854# 1.59e-20
C1803 xaa3.xa1b.MN0.D a_5844_56206# 0.0658f
C1804 AVDD xaa6.xg.XA7.MP1.G 2.06f
C1805 xaa6.xf.XA1.MN0.G xaa6.xg.XA4.MP0.D 3.2e-19
C1806 a_31132_56622# a_31132_56270# 0.0109f
C1807 a_37324_56622# xaa6.xg.XA6.MP0.D 0.00176f
C1808 xaa6.xd.XA7.MN1.D a_29764_55214# 0.00558f
C1809 xaa6.xd.XA1.MN0.G a_28612_55214# 1.17e-19
C1810 xaa3.xa1b.MN0.D a_4308_51566# 0.073f
C1811 PWRUP_1V8 xaa4.xa1.M3.D 6.23e-19
C1812 xaa6.xg.XA7.MN1.D xaa6.xg.XA4.MN0.D 0.026f
C1813 a_4692_56206# a_4692_55854# 0.0109f
C1814 AVDD a_26092_53806# 0.00164f
C1815 xaa1.xa4.M0.D m3_37668_110044# 0.074f
C1816 xaa6.xg.XA4.MN0.G xaa6.xg.XA3.MN1.G 0.0223f
C1817 xaa0.xa1.MN0.D xaa0.xa1.MP1.D 0.0657f
C1818 a_4692_58494# li_4980_58996# 2e-19
C1819 a_1220_74698# xaa1.xa3.D 0.00304f
C1820 a_n940_70022# a_788_72222# 2.35e-20
C1821 a_640_61158# xaa1.xb2.M7.D 0.00224f
C1822 a_n908_61510# xaa1.xa1.M1.D 6.46e-20
C1823 AVDD xaa3.xa4.MN0.D 0.72f
C1824 m2_4468_111644# m3_37748_111964# 0.0138f
C1825 PWRUP_1V8 xaa6.xf.XA4.MN0.D 0.00353f
C1826 xaa6.xg.XA7.MN1.G a_37324_56622# 0.0769f
C1827 xaa6.xg.XA7.MP1.G a_36172_56622# 0.0692f
C1828 xaa6.xd.XA1.MN0.G a_31132_56270# 0.00193f
C1829 a_36172_57326# a_36172_56974# 0.0109f
C1830 xaa6.xg.XA7.MN1.D xaa6.xg.XA6.MP0.D 0.0532f
C1831 xaa0.xa2a.MN0.D a_n908_53806# 1.31e-19
C1832 AVDD xaa6.xg.XA4.MN0.D 1.92e-19
C1833 xaa6.xf.XA5.MN0.G a_34804_55214# 0.0155f
C1834 xaa0.xa1.MN2.D a_n908_53806# 0.0472f
C1835 xaa0.xa1.MN0.D a_244_53806# 0.0889f
C1836 a_2948_70022# m1_4468_72124# 1.79e-19
C1837 xaa1.xa3.D m1_4468_71164# 12.9f
C1838 xaa1.xa4.M0.D m2_4468_105884# 71.5f
C1839 xaa1.xa4.M0.D m3_37748_76444# 0.111f
C1840 a_29764_53454# a_31132_53454# 8.89e-19
C1841 li_4468_84764# li_4468_84604# 7.91f
C1842 li_4468_109724# m1_4468_109724# 23f
C1843 xaa4.xa2.M0.G xaa5.xa3.xc1a.D 5.49e-20
C1844 xaa0.xa6.MN0.D xaa1.xa1.M3.D 8.17e-19
C1845 xaa3.xa1b.MN0.D xaa0.xa2a.MN0.D 0.00581f
C1846 CK a_29764_62510# 3.97e-20
C1847 xaa1.xa2.M5.D a_n908_61510# 8.62e-20
C1848 xaa1.xa2.M7.D PWRUP_1V8 2e-19
C1849 AVDD a_5844_63070# 0.388f
C1850 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MN1.G 0.311f
C1851 xaa6.xd.XA7.MN1.D a_29764_57326# 0.014f
C1852 PWRUP_1V8 xaa6.xf.XA6.MN0.D 0.00353f
C1853 xaa6.xf.XA1.MN0.G xaa6.xg.XA7.MP1.G 0.017f
C1854 a_31132_57678# xaa6.xe.XA7.MP1.G 2.36e-20
C1855 a_32284_57678# xaa6.xe.XA7.MN1.G 5.46e-19
C1856 AVDD xaa6.xg.XA6.MP0.D 0.147f
C1857 xaa6.xd.XA6.MN0.G xaa6.xd.XA5.MN0.G 0.27f
C1858 a_36172_56270# xaa6.xg.XA5.MN0.D 2.54e-19
C1859 xaa6.xg.XA7.MP1.G a_37324_54510# 0.0969f
C1860 xaa0.xa1.MN2.S a_244_53806# 0.00336f
C1861 xaa6.xd.XA1.MN0.G a_31132_53806# 0.00207f
C1862 xaa1.xa4.M0.D m3_4628_93564# 0.0276f
C1863 xaa1.xa4.M0.G xaa3.xa6.MN0.D 0.0148f
C1864 IBPSR_1U xaa3.xa1b.MN0.D 0.841f
C1865 xaa3.xa2.MN0.D xaa3.xa1capd.B 0.187f
C1866 a_4692_58142# a_5844_58142# 0.00133f
C1867 CK xaa6.xg.XA7.MN0.G 5.68e-19
C1868 PWRUP_1V8 xaa6.xf.XA7.MN1.G 0.667f
C1869 xaa3.xa1b.MN0.D a_4692_56206# 0.0782f
C1870 AVDD xaa6.xg.XA7.MN1.G 1.97f
C1871 m2_4468_98204# m3_37748_98524# 0.0138f
C1872 a_34804_57326# xaa6.xf.XA5.MN0.G 6.21e-20
C1873 xaa6.xf.XA1.MN0.G xaa6.xg.XA4.MN0.D 0.00287f
C1874 a_32284_56974# xaa6.xe.XA6.MN0.G 2.34e-19
C1875 xaa6.xd.XA7.MN1.D a_28612_55214# 0.00133f
C1876 xaa6.xc.XA1.MN0.G a_29764_55214# 1.02e-19
C1877 xaa1.xa4.M0.D li_4468_99004# 23f
C1878 IBPSR_1U a_4308_51566# 0.00731f
C1879 xaa3.xa1b.MN0.D a_4308_51918# 0.0751f
C1880 xaa6.xg.XA7.MN1.D xaa6.xg.XA4.MP1.G 0.00147f
C1881 a_4692_56206# a_5844_56206# 0.00133f
C1882 xaa1.xa4.M0.D m3_4788_110844# 0.0138f
C1883 a_29764_54862# xaa6.xd.XA3.MN0.D 0.00176f
C1884 a_36172_54862# a_37324_54862# 0.00133f
C1885 a_5844_58494# li_6204_59524# 1.49e-19
C1886 a_4692_58494# li_4836_58996# 4e-19
C1887 a_4308_51918# a_4308_51566# 0.0109f
C1888 a_n940_70022# a_356_70022# 9.03e-19
C1889 xaa1.xa1.M8.D xaa1.xa1.M2.D 0.0014f
C1890 m2_4468_111644# m3_37668_111964# 0.0138f
C1891 xaa6.xf.XA1.MN0.G xaa6.xg.XA6.MP0.D 3e-19
C1892 xaa6.xg.XA7.MN1.G a_36172_56622# 0.0111f
C1893 xaa6.xd.XA1.MN0.G a_29764_56270# 0.00204f
C1894 xaa6.xg.XA7.MN1.D xaa6.xg.XA6.MN0.D 0.0989f
C1895 xaa0.xa2a.MN0.D xaa0.xa1.MN2.D 1.67e-19
C1896 AVDD xaa6.xg.XA4.MP1.G 0.349f
C1897 xaa6.xf.XA5.MN0.G a_33652_55214# 0.00301f
C1898 xaa6.xf.XA6.MN0.G xaa6.xf.XA3.MP0.D 8.78e-20
C1899 xaa0.xa1.MN0.G a_n908_52750# 8.67e-19
C1900 xaa0.xa1.MN0.D a_n908_53806# 0.0715f
C1901 a_244_54158# a_244_53806# 0.0109f
C1902 a_34804_55566# xaa6.xf.XA4.MN0.D 0.00176f
C1903 a_27244_55566# a_27244_55214# 0.0109f
C1904 a_n908_54158# CK_REF 0.00164f
C1905 a_2948_70022# m1_4468_72284# 8.44e-19
C1906 xaa1.xa4.M0.D m2_4468_106844# 71.5f
C1907 xaa1.xa4.M0.D m3_37668_76444# 0.074f
C1908 a_27244_62862# xaa5.xa3.xb1_0.D 5.81e-19
C1909 xaa5.xa3.xb2_0.D a_27244_62510# 0.0683f
C1910 a_29764_62862# a_29764_62510# 0.0109f
C1911 IBPSR_1U xaa0.xa2a.MN0.D 0.58f
C1912 xaa5.xa3.xb1_0.G xaa5.xa3.xc1a.D 0.00129f
C1913 xaa5.xb1.MN1.G xaa5.xb1.MN0.D 0.0108f
C1914 AVDD a_4692_63070# 0.00171f
C1915 m1_4468_85724# m2_4468_85724# 12.9f
C1916 xaa6.xd.XA7.MN1.D a_28612_57326# 0.00337f
C1917 xaa6.xc.XA1.MN0.G a_29764_57326# 0.0662f
C1918 xaa6.xf.XA1.MN0.G xaa6.xg.XA7.MN1.G 0.128f
C1919 a_31132_57678# xaa6.xe.XA7.MN1.G 0.0736f
C1920 AVDD xaa6.xg.XA6.MN0.D 0.00913f
C1921 m2_4468_84764# m3_37748_85084# 0.0138f
C1922 xaa4.xa4.M0.D xaa4.xa1.M0.D 3.01e-19
C1923 a_32284_55918# a_33652_55918# 8.89e-19
C1924 xaa6.xd.XA7.MN1.G a_29764_54158# 0.0786f
C1925 xaa6.xg.XA7.MN1.G a_37324_54510# 0.00563f
C1926 xaa6.xg.XA7.MP1.G a_36172_54510# 0.0278f
C1927 xaa0.xa1.MN2.S a_n908_53806# 0.0398f
C1928 a_n908_55214# CK_REF 7.19e-20
C1929 xaa6.xd.XA1.MN0.G a_29764_53806# 0.0032f
C1930 a_34804_54158# a_36172_54158# 8.89e-19
C1931 xaa1.xa4.M0.D m3_37748_93724# 0.111f
C1932 li_4468_102044# li_4468_101884# 7.91f
C1933 xaa3.xa2.MN0.D a_5844_58142# 0.0897f
C1934 PWRUP_1V8 xaa6.xf.XA7.MP1.G 0.124f
C1935 IBPSR_1U a_4692_56206# 1.59e-20
C1936 AVDD xaa6.xf.XA7.MN0.D 0.486f
C1937 m2_4468_98204# m3_37668_98524# 0.0138f
C1938 xaa6.xf.XA1.MN0.G xaa6.xg.XA4.MP1.G 1.11e-19
C1939 a_29764_56622# a_29764_56270# 0.0109f
C1940 a_36172_56622# xaa6.xg.XA6.MN0.D 0.00176f
C1941 xaa6.xc.XA1.MN0.G a_28612_55214# 0.00196f
C1942 IBPSR_1U a_4308_51918# 0.136f
C1943 xaa3.xa1b.MN0.D xbb1.xa3.M0.D 1.38e-19
C1944 PWRUP_1V8 a_4308_53678# 1.25e-20
C1945 xaa6.xf.XA7.MN1.G a_34804_55566# 7.66e-19
C1946 AVDD xaa4.xa1.M3.D 0.00415f
C1947 xaa1.xa4.M0.D m3_4628_110844# 0.0276f
C1948 a_36172_55214# xaa6.xg.XA3.MN1.G 0.00114f
C1949 xaa0.xa2a.MN0.G a_n908_53102# 1.38e-19
C1950 xaa4.xa2.M0.D xaa4.xa1.M1.D 0.00147f
C1951 a_5844_58494# li_6132_59524# 4.95e-20
C1952 li_4468_87644# m1_4468_87644# 23f
C1953 xaa1.xa1.M5.D xaa0.xa2a.MN0.D 0.0105f
C1954 xaa5.xa3.xc1a.D a_27244_61102# 0.0467f
C1955 xaa1.xa1.M8.D xaa1.xb2.M0.D 0.0433f
C1956 AVDD xaa1.xb2.M0.D 0.0694f
C1957 xaa6.xf.XA1.MN0.G xaa6.xg.XA6.MN0.D 0.00272f
C1958 xaa6.xd.XA7.MN1.D a_29764_56270# 0.012f
C1959 xaa6.xd.XA1.MN0.G a_28612_56270# 1.17e-19
C1960 a_34804_57326# a_34804_56974# 0.0109f
C1961 xaa0.xa2a.MN0.D xaa0.xa1.MN0.D 0.00454f
C1962 AVDD xaa6.xf.XA4.MN0.D 1.92e-19
C1963 m2_4468_71324# m3_37748_71644# 0.0138f
C1964 xaa0.xa1.MN0.G a_244_53102# 0.0674f
C1965 xaa0.xa1.MN0.D xaa0.xa1.MN2.D 0.0093f
C1966 xaa1.xa3.D m1_4468_72124# 12.9f
C1967 xaa1.xa4.M0.D m2_4468_107804# 71.5f
C1968 xaa1.xa4.M0.D m3_4788_77244# 0.0138f
C1969 a_28612_53454# a_29764_53454# 0.00133f
C1970 xaa6.xg.XA1.MN0.D a_36172_53454# 0.0492f
C1971 xaa6.xc.XA1.MN0.D a_26092_53102# 0.00176f
C1972 li_4468_85564# li_4468_84764# 39.3f
C1973 a_26092_62862# xaa5.xa3.xb1_0.D 0.00139f
C1974 CK a_27244_62510# 0.00224f
C1975 xaa5.xa3.xb2_0.D a_26092_62510# 0.0972f
C1976 xaa1.xa2.M6.D a_n908_61510# 6.46e-20
C1977 xaa1.xa2.M7.D xaa1.xa1.M8.D 3.18e-19
C1978 IBPSR_1U xaa1.xa1.M5.D 0.026f
C1979 xaa0.xa6.MN0.D xaa1.xa1.M4.D 8.17e-19
C1980 xaa6.xc.XA1.MN0.G a_28612_57326# 0.0858f
C1981 xaa0.xa2a.MN0.D xaa0.xa1.MN2.S 0.0536f
C1982 xaa6.xf.XA7.MN1.D xaa6.xg.XA7.MN1.G 7.59e-20
C1983 IBPSR_1U xaa0.xa1.MN0.D 7.34e-20
C1984 xaa6.xg.XA7.MN1.D xaa6.xf.XA7.MN1.G 7.59e-20
C1985 AVDD xaa6.xf.XA6.MN0.D 0.00913f
C1986 m2_4468_84764# m3_37668_85084# 0.0138f
C1987 xaa6.xc.XA6.MN0.G xaa6.xc.XA5.MN0.G 0.27f
C1988 a_34804_56270# xaa6.xf.XA5.MN0.G 0.00131f
C1989 xaa6.xd.XA7.MP1.G a_29764_54158# 0.057f
C1990 xaa6.xd.XA7.MN1.G a_28612_54158# 0.0756f
C1991 xaa0.xa1.MN2.S xaa0.xa1.MN2.D 0.157f
C1992 xaa6.xd.XA7.MN1.D a_29764_53806# 3.97e-20
C1993 xaa6.xd.XA1.MN0.G a_28612_53806# 1.35e-19
C1994 xaa1.xa4.M0.D m3_37668_93724# 0.074f
C1995 xaa1.xa4.M0.G a_5844_63070# 1.28e-19
C1996 a_5844_63422# xaa3.xa1b.MN0.D 0.0658f
C1997 a_n908_63270# IBPSR_1U 0.0674f
C1998 a_5844_58494# a_5844_58142# 0.0109f
C1999 xaa3.xa2.MN0.D a_4692_58142# 0.117f
C2000 PWRUP_1V8 xaa6.xe.XA7.MN0.D 0.0493f
C2001 AVDD xaa6.xf.XA7.MN1.G 3.56f
C2002 xaa6.xf.XA1.MN0.G xaa6.xf.XA4.MN0.D 0.00303f
C2003 xaa6.xc.XA1.MN0.G a_27244_55214# 0.00207f
C2004 xaa1.xa4.M0.D li_4468_99964# 23f
C2005 IBPSR_1U xbb1.xa3.M0.D 0.0574f
C2006 xaa3.xa1b.MN0.D xbb1.xa3.M1.D 1.38e-19
C2007 PWRUP_1V8 a_244_52750# 4.63e-19
C2008 xaa6.xf.XA7.MP1.G a_34804_55566# 0.0964f
C2009 xaa6.xf.XA7.MN1.G a_33652_55566# 0.0769f
C2010 AVDD xaa4.xa1.M4.D 0.00415f
C2011 xaa1.xa4.M0.D m3_37748_111004# 0.111f
C2012 a_28612_54862# xaa6.xd.XA3.MP0.D 0.00176f
C2013 a_34804_54862# a_36172_54862# 8.89e-19
C2014 xbb1.xa3.M0.D a_4308_51918# 0.00155f
C2015 xaa1.xa4.M0.D a_788_72222# 2.72e-20
C2016 a_29764_61454# a_29764_61102# 0.0109f
C2017 PWRUP_1V8 xaa1.xa1.M3.D 5.67e-19
C2018 AVDD a_5844_60782# 0.348f
C2019 xaa6.xf.XA1.MN0.G xaa6.xf.XA6.MN0.D 0.00286f
C2020 PWRUP_1V8 xaa6.xe.XA4.MN0.D 0.00353f
C2021 xaa6.xf.XA7.MN0.D a_34804_56622# 1.28e-19
C2022 xaa6.xd.XA7.MN1.D a_28612_56270# 0.00378f
C2023 xaa6.xc.XA1.MN0.G a_29764_56270# 1.02e-19
C2024 xaa0.xa2a.MN0.D a_244_54158# 0.00172f
C2025 AVDD xaa6.xf.XA4.MP0.D 0.159f
C2026 m2_4468_71324# m3_37668_71644# 0.0138f
C2027 xaa6.xe.XA6.MN0.G xaa6.xe.XA3.MP0.D 8.78e-20
C2028 xaa6.xe.XA7.MN1.G a_32284_52750# 0.00154f
C2029 xaa0.xa1.MN0.G a_n908_53102# 0.0695f
C2030 a_n908_54158# a_n908_53806# 0.0109f
C2031 a_33652_55566# xaa6.xf.XA4.MP0.D 0.00176f
C2032 a_26092_55566# a_26092_55214# 0.0109f
C2033 a_n908_54510# CK_REF 7.36e-19
C2034 xaa1.xa3.D m1_4468_72284# 2.05e-19
C2035 xaa1.xa4.M0.D m2_4468_108764# 71.5f
C2036 xaa6.xe.XA5.MN0.G a_32284_55214# 0.00301f
C2037 xaa1.xa4.M0.D m3_4628_77244# 0.0276f
C2038 li_4468_110684# m1_4468_110684# 23f
C2039 CK a_26092_62510# 0.00357f
C2040 xaa5.xa3.xb2_0.D xaa5.xb2_2.MN0.D 0.00217f
C2041 a_28612_62862# a_28612_62510# 0.0109f
C2042 xaa5.xa3.xb2_0.G a_26092_61454# 0.074f
C2043 xaa4.xa2.M0.G a_29764_61454# 3.33e-19
C2044 AVDD xaa5.xb2_4.MN0.D 0.541f
C2045 m1_4468_86684# m2_4468_86684# 12.9f
C2046 PWRUP_1V8 xaa6.xe.XA6.MN0.D 0.00353f
C2047 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MN0.D 0.336f
C2048 a_29764_57678# xaa6.xd.XA7.MN0.D 0.00176f
C2049 xaa6.xf.XA1.MN0.G xaa6.xf.XA7.MN1.G 0.224f
C2050 xaa6.xc.XA1.MN0.G a_27244_57326# 0.00236f
C2051 xaa0.xa2a.MN0.D a_244_55214# 0.00301f
C2052 AVDD xaa6.xf.XA6.MP0.D 0.147f
C2053 a_11712_55918# xaa4.xa2.M0.D 0.0715f
C2054 a_31132_55918# a_32284_55918# 0.00133f
C2055 xaa6.xd.XA7.MP1.G a_28612_54158# 0.0545f
C2056 xaa6.xd.XA7.MN1.G a_27244_54158# 7.1e-20
C2057 xaa0.xa1.MN2.S xaa0.xa1.MN0.D 0.423f
C2058 xaa6.xd.XA7.MN1.D a_28612_53806# 0.0016f
C2059 xaa6.xc.XA1.MN0.G a_29764_53806# 1.11e-19
C2060 xaa6.xg.XA3.MN1.G a_37324_53806# 0.107f
C2061 a_33652_54158# a_34804_54158# 0.00133f
C2062 xaa1.xa4.M0.D m3_4788_94524# 0.0138f
C2063 li_4468_102844# li_4468_102044# 39.3f
C2064 xaa1.xa3.D xaa1.xa2.M3.D 0.00153f
C2065 xaa1.xa4.M0.G a_4692_63070# 0.00273f
C2066 a_4692_63422# xaa3.xa1b.MN0.D 0.0709f
C2067 PWRUP_1V8 xaa6.xe.XA7.MP1.G 0.124f
C2068 AVDD xaa6.xf.XA7.MP1.G 2.06f
C2069 xaa6.xf.XA1.MN0.G xaa6.xf.XA4.MP0.D 4.75e-19
C2070 xaa6.xf.XA7.MN1.D xaa6.xf.XA4.MN0.D 0.026f
C2071 a_28612_56622# a_28612_56270# 0.0109f
C2072 a_34804_56622# xaa6.xf.XA6.MN0.D 0.00176f
C2073 xaa6.xc.XA7.MN1.D a_27244_55214# 0.00133f
C2074 xaa6.xc.XA1.MN0.G a_26092_55214# 1.06e-19
C2075 IBPSR_1U xbb1.xa3.M1.D 0.0531f
C2076 xaa3.xa1b.MN0.D xbb1.xa3.M2.D 1.38e-19
C2077 PWRUP_1V8 a_n908_52750# 0.00163f
C2078 xaa6.xf.XA7.MP1.G a_33652_55566# 0.0292f
C2079 xaa6.xf.XA7.MN1.G a_32284_55566# 7.1e-20
C2080 AVDD a_4308_53678# 0.00227f
C2081 xaa1.xa4.M0.D m3_37668_111004# 0.074f
C2082 xaa0.xa2a.MN0.G a_n908_53454# 1.24e-19
C2083 a_37324_55918# m1_37504_55818# 0.0189f
C2084 xbb1.xa3.M1.D a_4308_51918# 5.84e-19
C2085 xaa1.xa4.M0.D a_356_70022# 6.05e-19
C2086 a_n940_70022# a_n76_72222# 0.00121f
C2087 a_n908_61510# xaa1.xa1.M2.D 8.62e-20
C2088 AVDD a_4692_60782# 0.00171f
C2089 xaa6.xf.XA1.MN0.G xaa6.xf.XA6.MP0.D 4.47e-19
C2090 PWRUP_1V8 xaa6.xd.XA4.MN0.D 0.00353f
C2091 xaa6.xf.XA7.MN1.D xaa6.xf.XA6.MN0.D 0.0989f
C2092 xaa4.xa4.M0.D xaa4.xa2.M0.D 1.68f
C2093 xaa6.xf.XA7.MN0.D a_33652_56622# 0.0217f
C2094 xaa6.xf.XA7.MN1.G a_34804_56622# 0.0111f
C2095 xaa6.xc.XA1.MN0.G a_28612_56270# 0.00211f
C2096 a_33652_57326# a_33652_56974# 0.0109f
C2097 xaa0.xa2a.MN0.D a_n908_54158# 2.92e-19
C2098 AVDD xaa6.xe.XA4.MP0.D 0.159f
C2099 xaa6.xe.XA7.MN1.G a_31132_52750# 2.64e-19
C2100 xaa0.xa1.MN0.G a_244_53454# 0.066f
C2101 a_244_54158# xaa0.xa1.MN0.D 0.0658f
C2102 a_n908_54158# xaa0.xa1.MN2.D 0.00176f
C2103 xaa0.xa2a.MN0.G CK_REF 0.00875f
C2104 xaa1.xa4.M0.D m2_4468_109724# 71.5f
C2105 xaa6.xe.XA5.MN0.G a_31132_55214# 0.0155f
C2106 xaa1.xa4.M0.D m3_37748_77404# 0.111f
C2107 a_27244_53454# a_28612_53454# 8.89e-19
C2108 xaa6.xf.XA1.MN0.D a_34804_53454# 0.0492f
C2109 xaa6.xg.XA7.MN0.G m1_37504_55818# 6.41e-20
C2110 li_4468_85724# li_4468_85564# 7.91f
C2111 CK xaa5.xb2_2.MN0.D 7.29e-20
C2112 xaa1.xa3.D xaa1.xb1.M0.D 1.22e-19
C2113 xaa4.xa2.M0.G a_28612_61454# 0.0543f
C2114 AVDD a_29764_63566# 0.00139f
C2115 PWRUP_1V8 xaa6.xd.XA6.MN0.D 0.00353f
C2116 xaa6.xc.XA1.MN0.G a_26092_57326# 1.06e-19
C2117 a_28612_57678# xaa6.xd.XA7.MN0.D 0.00176f
C2118 a_29764_57678# xaa6.xd.XA7.MN1.G 0.072f
C2119 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MN1.G 0.467f
C2120 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN0.D 0.129f
C2121 xaa6.xf.XA1.MN0.G xaa6.xf.XA7.MP1.G 0.0184f
C2122 xaa6.xc.XA7.MN1.D a_27244_57326# 0.00337f
C2123 xaa0.xa5.MN2.G a_28612_57326# 2.93e-19
C2124 xaa0.xa2a.MN0.D a_n908_55214# 3.72e-19
C2125 AVDD xaa6.xe.XA6.MP0.D 0.147f
C2126 xaa0.xa1.MN2.S a_244_54158# 0.0893f
C2127 xaa6.xc.XA1.MN0.G a_28612_53806# 0.00209f
C2128 xaa6.xg.XA3.MN1.G a_36172_53806# 0.113f
C2129 a_10092_54510# xaa4.xa1.M1.D 6.46e-20
C2130 xaa1.xa4.M0.D m3_4628_94524# 0.0276f
C2131 a_5844_58494# xaa3.xa2.MN0.D 0.0658f
C2132 a_4692_58494# a_4692_58142# 0.0109f
C2133 PWRUP_1V8 xaa6.xe.XA7.MN1.G 0.658f
C2134 AVDD xaa6.xe.XA7.MN0.D 0.485f
C2135 xaa6.xe.XA1.MN0.G xaa6.xf.XA4.MN0.D 3.2e-19
C2136 xaa6.xf.XA7.MN1.D xaa6.xf.XA4.MP0.D 0.00426f
C2137 a_28612_56974# xaa6.xd.XA6.MN0.G 2.34e-19
C2138 xaa6.xc.XA7.MN1.D a_26092_55214# 0.00558f
C2139 xaa1.xa4.M0.D li_4468_100924# 23f
C2140 IBPSR_1U xbb1.xa3.M2.D 0.0506f
C2141 a_31132_57326# xaa6.xe.XA5.MN0.G 6.98e-20
C2142 a_244_55214# xaa0.xa1.MN2.S 0.0658f
C2143 AVDD a_244_52750# 0.443f
C2144 xaa1.xa4.M0.D m3_4788_111804# 0.0138f
C2145 a_27244_54862# xaa6.xc.XA3.MP0.D 0.00176f
C2146 a_33652_54862# a_34804_54862# 0.00133f
C2147 xbb1.xa3.M2.D a_4308_51918# 2.99e-19
C2148 xbb1.xa3.M1.D xbb1.xa3.M0.D 0.0488f
C2149 a_n940_70022# a_n508_70022# 0.00813f
C2150 li_4468_88604# m1_4468_88604# 23f
C2151 a_640_61158# xaa0.xa2a.MN0.D 0.0725f
C2152 a_28612_61454# a_28612_61102# 0.0109f
C2153 xaa1.xa1.M8.D xaa1.xa1.M3.D 0.00177f
C2154 PWRUP_1V8 xaa1.xa1.M4.D 5.67e-19
C2155 m2_4468_112604# m3_37748_112924# 0.0138f
C2156 xaa6.xe.XA1.MN0.G xaa6.xf.XA6.MN0.D 3e-19
C2157 xaa6.xf.XA7.MN1.D xaa6.xf.XA6.MP0.D 0.0532f
C2158 xaa6.xf.XA7.MN1.G a_33652_56622# 0.0785f
C2159 xaa6.xf.XA7.MP1.G a_34804_56622# 0.0676f
C2160 xaa6.xc.XA1.MN0.G a_27244_56270# 0.00207f
C2161 xaa0.xa2a.MN0.D a_244_54510# 0.00581f
C2162 AVDD xaa6.xe.XA4.MN0.D 1.92e-19
C2163 xaa0.xa1.MN0.G a_n908_53454# 0.0676f
C2164 xaa4.xa1.M8.D a_10092_55038# 0.0548f
C2165 a_n908_54158# xaa0.xa1.MN0.D 0.0675f
C2166 a_32284_55566# xaa6.xe.XA4.MP0.D 0.00176f
C2167 xaa1.xa4.M0.D m2_4468_110684# 71.5f
C2168 xaa1.xa4.M0.D m3_37668_77404# 0.074f
C2169 xaa4.xa1.M3.D a_10092_52750# 1.81e-19
C2170 xaa6.xg.XA7.MN0.G m1_37504_57930# 0.0488f
C2171 xaa5.xb2_3.MN0.D a_29764_62510# 0.00263f
C2172 a_29764_62862# xaa5.xb2_2.MN0.D 0.0682f
C2173 a_27244_62862# a_27244_62510# 0.0109f
C2174 xaa4.xa2.M0.G a_27244_61454# 5.56e-19
C2175 xaa1.xa2.M7.D a_n908_61510# 5.02e-20
C2176 CK xaa5.xa3.xb2_0.D 0.0746f
C2177 xaa5.xb1.MN1.G a_29764_61454# 0.0766f
C2178 IBPSR_1U a_640_61158# 6.96e-19
C2179 AVDD a_28612_63566# 0.351f
C2180 m1_4468_87644# m2_4468_87644# 12.9f
C2181 a_28612_57678# xaa6.xd.XA7.MN1.G 5.46e-19
C2182 a_29764_57678# xaa6.xd.XA7.MP1.G 2.36e-20
C2183 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MP1.G 0.313f
C2184 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN1.G 0.201f
C2185 xaa0.xa5.MN2.G a_27244_57326# 0.081f
C2186 xaa6.xc.XA7.MN1.D a_26092_57326# 0.014f
C2187 a_36172_57678# a_37324_57678# 0.00133f
C2188 xaa0.xa2a.MN0.D xaa0.xa3.MP0.D 5.08e-19
C2189 AVDD xaa6.xe.XA6.MN0.D 0.00913f
C2190 xaa6.xf.XA7.MN1.G a_34804_54510# 0.0835f
C2191 a_29764_55918# a_31132_55918# 8.89e-19
C2192 xaa6.xg.XA6.MN0.G a_37324_55918# 0.0674f
C2193 xaa0.xa1.MN2.S a_n908_54158# 0.0974f
C2194 xaa6.xc.XA1.MN0.G a_27244_53806# 0.0044f
C2195 xaa0.xa1.MN0.G CK_REF 0.13f
C2196 a_32284_54158# a_33652_54158# 8.89e-19
C2197 xaa1.xa4.M0.D m3_37748_94684# 0.111f
C2198 li_4468_103004# li_4468_102844# 7.91f
C2199 xaa1.xa2.M8.D IBPSR_1U 0.0166f
C2200 xaa3.xa8.MP0.D xaa3.xa1b.MN0.D 0.00994f
C2201 xaa1.xa3.D xaa1.xa2.M4.D 0.00203f
C2202 PWRUP_1V8 xaa6.xd.XA7.MN0.D 0.0493f
C2203 a_4692_58494# xaa3.xa2.MN0.D 0.0728f
C2204 AVDD xaa6.xe.XA7.MP1.G 2.06f
C2205 m2_4468_99164# m3_37748_99484# 0.0138f
C2206 xaa6.xe.XA1.MN0.G xaa6.xf.XA4.MP0.D 0.00287f
C2207 a_27244_56622# a_27244_56270# 0.0109f
C2208 a_33652_56622# xaa6.xf.XA6.MP0.D 0.00176f
C2209 PWRUP_1V8 a_n908_53102# 0.00117f
C2210 a_n908_55214# xaa0.xa1.MN2.S 0.0702f
C2211 AVDD a_n908_52750# 0.00527f
C2212 xaa1.xa4.M0.D m3_4628_111804# 0.0276f
C2213 xaa1.xa1.M6.D xaa0.xa2a.MN0.D 0.0116f
C2214 xaa1.xa1.M8.D a_640_60806# 0.0871f
C2215 AVDD a_640_60806# 0.356f
C2216 m2_4468_112604# m3_37668_112924# 0.0138f
C2217 xaa6.xe.XA1.MN0.G xaa6.xf.XA6.MP0.D 0.00276f
C2218 xaa6.xc.XA7.MN1.D a_27244_56270# 0.00378f
C2219 xaa6.xf.XA7.MP1.G a_33652_56622# 0.029f
C2220 xaa6.xc.XA1.MN0.G a_26092_56270# 1.06e-19
C2221 a_n908_56270# a_244_56270# 0.00133f
C2222 a_32284_57326# a_32284_56974# 0.0109f
C2223 xaa0.xa2a.MN0.D a_n908_54510# 0.00305f
C2224 AVDD xaa6.xd.XA4.MN0.D 1.92e-19
C2225 xaa6.xg.XA7.MP1.G a_36172_53102# 1.1e-19
C2226 xaa6.xg.XA7.MN1.G a_37324_53102# 0.00531f
C2227 xaa0.xa1.MN0.G xaa0.xa1.MP1.D 0.0106f
C2228 a_n908_54158# a_244_54158# 0.00133f
C2229 xaa0.xa2a.MN0.G a_n908_53806# 8.26e-19
C2230 a_n908_54862# CK_REF 2.53e-19
C2231 xaa1.xa4.M0.D m2_4468_111644# 71.5f
C2232 xaa6.xd.XA5.MN0.G a_29764_55214# 0.0155f
C2233 xaa1.xa4.M0.D m3_4788_78204# 0.0138f
C2234 a_26092_53454# a_27244_53454# 0.00133f
C2235 xaa4.xa1.M4.D a_10092_52750# 1.21e-19
C2236 li_4468_86524# li_4468_85724# 39.3f
C2237 li_4468_111644# m1_4468_111644# 23f
C2238 a_27244_63214# xaa5.xa3.xb1_0.D 2.74e-19
C2239 xaa5.xb2_3.MN0.D a_28612_62510# 0.00224f
C2240 a_28612_62862# xaa5.xb2_2.MN0.D 0.0674f
C2241 xaa5.xa3.xb1_0.G a_27244_61454# 3.13e-19
C2242 xaa5.xb1.MN1.G a_28612_61454# 0.0684f
C2243 IBPSR_1U xaa1.xa1.M6.D 0.026f
C2244 AVDD xaa5.xa3.xb2_0.G 0.952f
C2245 a_28612_57678# xaa6.xd.XA7.MP1.G 0.071f
C2246 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MP1.G 0.216f
C2247 xaa6.xe.XA7.MN1.D xaa6.xf.XA7.MN1.G 1.74e-19
C2248 xaa0.xa5.MN2.G a_26092_57326# 0.0678f
C2249 xaa0.xa2a.MN0.D a_244_55566# 0.00147f
C2250 AVDD xaa6.xd.XA6.MN0.D 0.00913f
C2251 m2_4468_85724# m3_37748_86044# 0.0138f
C2252 xaa6.xf.XA7.MN1.G a_33652_54510# 0.0057f
C2253 xaa6.xf.XA7.MP1.G a_34804_54510# 0.0278f
C2254 xaa6.xc.XA7.MP1.G a_27244_54158# 0.0545f
C2255 xaa6.xc.XA7.MN1.G a_28612_54158# 7.1e-20
C2256 a_31132_56270# xaa6.xe.XA5.MN0.G 0.00131f
C2257 xaa6.xc.XA7.MN1.D a_27244_53806# 0.0016f
C2258 xaa6.xg.XA6.MN0.G a_36172_55918# 0.0658f
C2259 xaa0.xa1.MN2.S a_244_54510# 0.0662f
C2260 xaa6.xc.XA1.MN0.G a_26092_53806# 0.00318f
C2261 xaa0.xa1.MN0.G a_244_53806# 2.33e-19
C2262 xaa1.xa4.M0.D m3_37668_94684# 0.074f
C2263 a_37324_54862# m1_37504_55818# 0.00375f
C2264 xaa3.xa7.MN0.D xaa3.xa1b.MN0.D 0.123f
C2265 a_4692_63422# a_5844_63422# 0.00133f
C2266 xaa1.xa2.M8.D a_n908_63270# 0.0534f
C2267 PWRUP_1V8 xaa6.xd.XA7.MN1.G 0.667f
C2268 a_4692_58494# a_5844_58494# 0.00133f
C2269 AVDD xaa6.xe.XA7.MN1.G 3.52f
C2270 m2_4468_99164# m3_37668_99484# 0.0138f
C2271 xaa6.xe.XA7.MN1.G a_33652_55566# 7.1e-20
C2272 xaa6.xe.XA7.MP1.G a_32284_55566# 0.0292f
C2273 xaa1.xa4.M0.D li_4468_101884# 23f
C2274 xaa4.xa4.M0.D a_10092_54510# 1.74e-19
C2275 a_29764_57326# xaa6.xd.XA5.MN0.G 6.21e-20
C2276 a_n908_55214# a_244_55214# 0.00133f
C2277 xaa0.xa3.MP0.D xaa0.xa1.MN2.S 0.00987f
C2278 a_27244_56974# xaa6.xc.XA6.MN0.G 2.34e-19
C2279 xaa6.xe.XA1.MN0.G xaa6.xe.XA4.MP0.D 0.00303f
C2280 AVDD a_244_53102# 0.485f
C2281 xaa1.xa4.M0.D m3_37748_111964# 0.111f
C2282 a_26092_54862# xaa6.xc.XA3.MN0.D 0.00176f
C2283 a_32284_54862# a_33652_54862# 8.89e-19
C2284 xbb1.xa3.M2.D xbb1.xa3.M1.D 0.0488f
C2285 xaa1.xa4.M0.D a_n76_72222# 0.00214f
C2286 xaa1.xa1.M6.D xaa1.xa1.M5.D 0.0488f
C2287 xaa5.xa3.xb1_0.D a_27244_60750# 0.00102f
C2288 PWRUP_1V8 a_29764_61102# 0.0699f
C2289 a_27244_61454# a_27244_61102# 0.0109f
C2290 xaa1.xa1.M8.D xaa1.xa1.M4.D 0.00232f
C2291 xaa6.xe.XA1.MN0.G xaa6.xe.XA6.MP0.D 0.00286f
C2292 PWRUP_1V8 xaa6.xc.XA4.MN0.D 0.00353f
C2293 xaa0.xa5.MN2.G a_27244_56270# 1.49e-19
C2294 xaa6.xc.XA7.MN1.D a_26092_56270# 0.012f
C2295 xaa0.xa2a.MN0.D xaa0.xa2a.MN0.G 0.14f
C2296 AVDD xaa6.xd.XA4.MP0.D 0.159f
C2297 m2_4468_72284# m3_37748_72604# 0.0138f
C2298 xaa6.xd.XA6.MN0.G xaa6.xd.XA3.MP0.D 8.78e-20
C2299 xaa6.xd.XA7.MN1.G a_29764_52750# 2.64e-19
C2300 a_244_54510# a_244_54158# 0.0109f
C2301 a_31132_55566# xaa6.xe.XA4.MN0.D 0.00176f
C2302 xaa6.xg.XA5.MN0.G xaa6.xg.XA4.MP0.D 0.0618f
C2303 xaa1.xa4.M0.D m2_4468_112604# 71.5f
C2304 xaa6.xd.XA5.MN0.G a_28612_55214# 0.00301f
C2305 xaa1.xa4.M0.D m3_4628_78204# 0.0276f
C2306 a_26092_63214# xaa5.xa3.xb1_0.D 5.31e-19
C2307 a_26092_62862# a_26092_62510# 0.0109f
C2308 xaa5.xa3.xb1_0.G a_26092_61454# 0.0752f
C2309 xaa4.xa2.M0.G PWRUP_1V8 0.0305f
C2310 xaa1.xa3.D a_640_60278# 5.46e-19
C2311 a_29764_62862# CK 3.97e-20
C2312 AVDD a_29764_63918# 0.00139f
C2313 m1_4468_88604# m2_4468_88604# 12.9f
C2314 PWRUP_1V8 xaa6.xc.XA6.MN0.D 0.00353f
C2315 xaa6.xe.XA1.MN0.G xaa6.xe.XA7.MN0.D 0.00664f
C2316 xaa0.xa2a.MN0.D a_n908_55566# 2.13e-19
C2317 a_34804_57678# a_36172_57678# 8.89e-19
C2318 AVDD xaa6.xd.XA6.MP0.D 0.147f
C2319 m2_4468_85724# m3_37668_86044# 0.0138f
C2320 xaa6.xf.XA7.MP1.G a_33652_54510# 0.0953f
C2321 xaa6.xf.XA7.MN1.G a_32284_54510# 7.1e-20
C2322 xaa6.xc.XA7.MP1.G a_26092_54158# 0.057f
C2323 xaa6.xc.XA7.MN1.G a_27244_54158# 0.074f
C2324 xaa6.xc.XA7.MN1.D a_26092_53806# 3.97e-20
C2325 xaa0.xa1.MN2.S a_n908_54510# 0.0978f
C2326 xaa0.xa1.MN0.G a_n908_53806# 0.00507f
C2327 a_28612_55918# a_29764_55918# 0.00133f
C2328 a_31132_54158# a_32284_54158# 0.00133f
C2329 xaa1.xa4.M0.D m3_4788_95484# 0.0138f
C2330 li_4468_103804# li_4468_103004# 39.3f
C2331 PWRUP_1V8 xaa6.xd.XA7.MP1.G 0.124f
C2332 AVDD xaa6.xd.XA7.MN0.D 0.485f
C2333 xaa6.xe.XA7.MP1.G a_31132_55566# 0.098f
C2334 xaa6.xe.XA7.MN1.G a_32284_55566# 0.0754f
C2335 xaa6.xg.XA7.MP1.G xaa6.xg.XA5.MN0.G 0.397f
C2336 xaa0.xa3.MP0.D a_244_55214# 0.0494f
C2337 a_32284_56622# xaa6.xe.XA6.MP0.D 0.00176f
C2338 a_26092_56622# a_26092_56270# 0.0109f
C2339 xaa6.xe.XA7.MN1.D xaa6.xe.XA4.MP0.D 0.00426f
C2340 xaa6.xe.XA1.MN0.G xaa6.xe.XA4.MN0.D 4.75e-19
C2341 AVDD a_n908_53102# 0.00171f
C2342 xaa1.xa4.M0.D m3_37668_111964# 0.074f
C2343 xaa1.xa4.M0.D a_n508_70022# 0.00673f
C2344 li_4468_89564# m1_4468_89564# 23f
C2345 xaa5.xa3.xb1_0.D a_26092_60750# 0.00404f
C2346 xaa1.xa1.M8.D xaa1.xb2.M7.D 0.043f
C2347 PWRUP_1V8 a_28612_61102# 0.0674f
C2348 a_n908_61510# xaa1.xa1.M3.D 1.21e-19
C2349 AVDD xaa1.xb2.M7.D 0.166f
C2350 xaa6.xe.XA1.MN0.G xaa6.xe.XA6.MN0.D 4.47e-19
C2351 xaa6.xe.XA7.MN1.D xaa6.xe.XA6.MP0.D 0.0532f
C2352 PWRUP_1V8 CK_REF 0.0418f
C2353 xaa4.xa2.M0.G a_11712_54334# 0.00555f
C2354 xaa6.xg.XA7.MN0.D a_37324_56974# 0.016f
C2355 xaa0.xa5.MN2.D a_n908_56270# 0.0492f
C2356 xaa0.xa5.MN0.D a_244_56270# 0.0889f
C2357 a_31132_57326# a_31132_56974# 0.0109f
C2358 xaa0.xa2a.MN0.D a_244_54862# 0.0297f
C2359 xaa6.xe.XA7.MN0.D a_32284_56622# 0.0217f
C2360 AVDD xaa6.xc.XA4.MP0.D 0.159f
C2361 m2_4468_72284# m3_37668_72604# 0.0138f
C2362 xaa0.xa2a.MN0.G xaa0.xa1.MN0.D 0.00197f
C2363 xaa6.xg.XA5.MN0.G xaa6.xg.XA4.MN0.D 0.126f
C2364 xaa1.xa4.M0.D m2_4468_113564# 71.5f
C2365 xaa6.xd.XA7.MN1.G a_28612_52750# 0.00154f
C2366 xaa1.xa4.M0.D m3_37748_78364# 0.111f
C2367 a_4308_53678# xbb1.xa3.M3.D 1.21e-19
C2368 a_37324_53806# a_37324_53454# 0.0109f
C2369 xaa6.xe.XA1.MN0.D a_31132_53454# 0.0492f
C2370 li_4468_86684# li_4468_86524# 7.91f
C2371 xaa0.xa6.MN0.D xaa0.xa2a.MN0.D 3.25f
C2372 xaa1.xa2.M3.D xaa1.xa2.M2.D 0.0488f
C2373 a_27244_62862# xaa5.xa3.xb2_0.D 0.066f
C2374 AVDD a_28612_63918# 0.351f
C2375 PWRUP_1V8 a_5844_55854# 0.0658f
C2376 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MN0.D 0.336f
C2377 a_27244_57678# xaa6.xc.XA7.MN0.D 0.00176f
C2378 xaa0.xa2a.MN0.D xaa0.xa1.MN0.G 0.0446f
C2379 xaa6.xd.XA1.MN0.G xaa6.xf.XA7.MP1.G 4.23e-19
C2380 xaa6.xf.XA7.MN1.D xaa6.xe.XA7.MN1.G 1.74e-19
C2381 xaa6.xe.XA1.MN0.G xaa6.xe.XA7.MP1.G 0.027f
C2382 AVDD xaa6.xc.XA6.MP0.D 0.147f
C2383 xaa6.xc.XA7.MN1.G a_26092_54158# 0.0802f
C2384 xaa6.xf.XA6.MN0.G a_34804_55918# 0.0889f
C2385 xaa0.xa1.MN2.S xaa0.xa2a.MN0.G 0.405f
C2386 xaa0.xa1.MN0.G xaa0.xa1.MN2.D 0.00321f
C2387 a_29764_56270# xaa6.xd.XA5.MN0.G 0.00131f
C2388 xaa1.xa4.M0.D m3_4628_95484# 0.0276f
C2389 xaa0.xa6.MN0.D IBPSR_1U 0.226f
C2390 xaa3.xa8.MP0.D a_5844_63422# 0.0494f
C2391 xaa1.xa3.D xaa1.xa2.M5.D 0.00279f
C2392 PWRUP_1V8 xaa6.xc.XA7.MN0.D 0.0497f
C2393 IBPSR_1U xaa0.xa1.MN0.G 0.00162f
C2394 AVDD xaa6.xd.XA7.MN1.G 3.56f
C2395 xaa6.xe.XA7.MN1.G a_31132_55566# 7.66e-19
C2396 xaa6.xd.XA1.MN0.G xaa6.xe.XA4.MP0.D 3.2e-19
C2397 a_n908_55566# xaa0.xa1.MN2.S 2.92e-19
C2398 xaa1.xa4.M0.D li_4468_102844# 23f
C2399 xaa6.xg.XA7.MP1.G xaa6.xg.XA5.MN0.D 0.0398f
C2400 a_244_55566# a_244_55214# 0.0109f
C2401 xaa6.xe.XA7.MN1.D xaa6.xe.XA4.MN0.D 0.026f
C2402 xaa6.xg.XA7.MN1.G xaa6.xg.XA5.MN0.G 0.0247f
C2403 AVDD a_244_53454# 0.365f
C2404 xaa1.xa4.M0.D m3_4788_112764# 0.0138f
C2405 xaa4.xa2.M0.D xaa4.xa1.M2.D 0.00187f
C2406 a_31132_54862# a_32284_54862# 0.00133f
C2407 li_4468_70204# li_4468_69404# 39.3f
C2408 a_29764_61454# xaa5.xb1.MN0.D 0.00176f
C2409 a_26092_61454# a_26092_61102# 0.0109f
C2410 AVDD a_29764_61102# 0.00132f
C2411 xaa6.xg.XA7.MP1.G a_37324_56974# 0.0291f
C2412 xaa6.xe.XA7.MN1.D xaa6.xe.XA6.MN0.D 0.0989f
C2413 xaa6.xd.XA1.MN0.G xaa6.xe.XA6.MP0.D 3.43e-19
C2414 xaa6.xe.XA7.MP1.G a_32284_56622# 0.029f
C2415 xaa6.xg.XA7.MN0.D a_36172_56974# 0.00297f
C2416 xaa0.xa5.MN0.D a_n908_56270# 0.073f
C2417 a_244_56622# a_244_56270# 0.0109f
C2418 a_37324_57326# xaa6.xg.XA7.MN0.G 0.0658f
C2419 a_36172_57326# xaa6.xg.XA7.MN2.D 0.00176f
C2420 xaa0.xa2a.MN0.D a_n908_54862# 0.0297f
C2421 xaa6.xe.XA7.MN0.D a_31132_56622# 1.28e-19
C2422 AVDD xaa6.xc.XA4.MN0.D 1.92e-19
C2423 xaa6.xc.XA6.MN0.G xaa6.xc.XA3.MP0.D 8.78e-20
C2424 xaa6.xg.XA5.MN0.G xaa6.xg.XA4.MP1.G 0.034f
C2425 xaa0.xa2a.MN0.G a_244_54158# 0.00224f
C2426 a_n908_54510# a_n908_54158# 0.0109f
C2427 a_29764_55566# xaa6.xd.XA4.MN0.D 0.00176f
C2428 xaa1.xa4.M0.D m2_4468_114524# 71.5f
C2429 xaa6.xc.XA5.MN0.G a_27244_55214# 0.00301f
C2430 xaa1.xa4.M0.D m3_37668_78364# 0.074f
C2431 li_4468_112604# m1_4468_112604# 23f
C2432 xaa5.xb2_3.MN0.D xaa5.xb2_2.MN0.D 0.197f
C2433 xaa5.xb1.MN1.G PWRUP_1V8 0.088f
C2434 xaa0.xa6.MN0.D xaa1.xa1.M5.D 7.41e-19
C2435 a_26092_62862# xaa5.xa3.xb2_0.D 0.0711f
C2436 a_27244_62862# CK 0.0234f
C2437 a_28612_62862# a_29764_62862# 0.00133f
C2438 AVDD xaa4.xa2.M0.G 10.3f
C2439 m1_4468_89564# m2_4468_89564# 12.9f
C2440 PWRUP_1V8 a_4692_55854# 0.0674f
C2441 a_26092_57678# xaa6.xc.XA7.MN0.D 0.00176f
C2442 xaa0.xa2a.MN0.D a_244_55918# 9.04e-19
C2443 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN0.D 0.12f
C2444 a_37324_58030# xaa6.xg.XA7.MP1.G 3.8e-19
C2445 xaa1.xa3.D a_10092_55038# 0.0705f
C2446 xaa6.xe.XA1.MN0.G xaa6.xe.XA7.MN1.G 0.412f
C2447 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MP1.G 0.313f
C2448 a_33652_57678# a_34804_57678# 0.00133f
C2449 a_27244_57678# xaa6.xc.XA7.MP1.G 0.0694f
C2450 AVDD xaa6.xc.XA6.MN0.D 0.00913f
C2451 xaa6.xf.XA6.MN0.G a_33652_55918# 0.111f
C2452 xaa0.xa1.MN2.S a_244_54862# 0.0678f
C2453 xaa0.xa1.MN0.G xaa0.xa1.MN0.D 0.274f
C2454 a_27244_55918# a_28612_55918# 8.89e-19
C2455 a_29764_54158# a_31132_54158# 8.89e-19
C2456 xaa1.xa4.M0.D m3_37748_95644# 0.111f
C2457 li_4468_103964# li_4468_103804# 7.91f
C2458 xaa0.xa6.MN0.D a_n908_63270# 0.0714f
C2459 xaa3.xa7.MN0.D a_5844_63422# 0.0677f
C2460 xaa5.xb3.MP1.D xaa5.xb2_4.MN0.D 1.42e-19
C2461 PWRUP_1V8 xaa6.xc.XA7.MP1.G 0.124f
C2462 AVDD xaa6.xd.XA7.MP1.G 2.06f
C2463 xaa6.xd.XA1.MN0.G xaa6.xe.XA4.MN0.D 0.00287f
C2464 xaa6.xg.XA7.MN1.G xaa6.xg.XA5.MN0.D 0.00451f
C2465 CK xaa6.xg.XA1.MN0.D 0.0112f
C2466 xaa0.xa1.MN0.G xaa0.xa1.MN2.S 0.094f
C2467 a_31132_56622# xaa6.xe.XA6.MN0.D 0.00176f
C2468 AVDD a_n908_53454# 0.00164f
C2469 xaa6.xg.XA4.MN0.G a_37324_54862# 0.0674f
C2470 xaa1.xa4.M0.D m3_4628_112764# 0.0276f
C2471 xaa1.xa4.M0.D a_n940_70022# 0.181f
C2472 xaa5.xb1.MN1.D a_29764_61102# 0.0126f
C2473 a_n908_61510# xaa1.xa1.M4.D 1.81e-19
C2474 AVDD a_28612_61102# 0.352f
C2475 m2_4468_113564# m3_37748_113884# 0.0138f
C2476 xaa6.xg.XA7.MN1.G a_37324_56974# 0.0035f
C2477 xaa6.xg.XA7.MP1.G a_36172_56974# 2.35e-19
C2478 IBPSR_1U xaa4.xa1.M5.D 0.026f
C2479 xaa6.xd.XA1.MN0.G xaa6.xe.XA6.MN0.D 0.00272f
C2480 xaa6.xe.XA7.MN1.G a_32284_56622# 0.0769f
C2481 xaa6.xe.XA7.MP1.G a_31132_56622# 0.0692f
C2482 a_36172_57326# xaa6.xg.XA7.MN0.G 0.0674f
C2483 a_29764_57326# a_29764_56974# 0.0109f
C2484 xaa0.xa5.MN0.D xaa0.xa5.MN2.D 0.0215f
C2485 AVDD CK_REF 0.562f
C2486 xaa0.xa2a.MN0.G a_n908_54158# 0.00459f
C2487 a_n908_54510# a_244_54510# 0.00133f
C2488 xaa1.xa4.M0.D m2_4468_115484# 71.5f
C2489 xaa6.xf.XA7.MN1.G a_34804_53102# 7.28e-19
C2490 xaa6.xc.XA5.MN0.G a_26092_55214# 0.0155f
C2491 xaa6.xd.XA1.MN0.D a_29764_53454# 0.0492f
C2492 a_36172_53806# a_36172_53454# 0.0109f
C2493 xaa1.xa4.M0.D m3_4788_79164# 0.0138f
C2494 li_4468_87484# li_4468_86684# 39.3f
C2495 xaa4.xa2.M0.G xaa5.xb1.MN1.D 0.226f
C2496 xaa3.xa1b.MN0.D PWRUP_1V8 1.73f
C2497 a_26092_62862# CK 0.0374f
C2498 AVDD xaa5.xa3.xb1_0.G 0.826f
C2499 xaa0.xa2a.MN0.D a_n908_55918# 1.17e-19
C2500 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MP1.G 0.21f
C2501 a_37324_58030# xaa6.xg.XA7.MN1.G 4.26e-19
C2502 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MN1.G 0.467f
C2503 a_26092_57678# xaa6.xc.XA7.MP1.G 2.36e-20
C2504 a_27244_57678# xaa6.xc.XA7.MN1.G 5.46e-19
C2505 AVDD a_5844_55854# 0.388f
C2506 PWRUP_1V8 a_4308_51566# 0.0105f
C2507 xaa6.xg.XA7.MP1.G xaa6.xg.XA3.MP0.D 0.0712f
C2508 a_37324_56270# a_37324_55918# 0.0109f
C2509 xaa0.xa1.MN2.S a_n908_54862# 0.0962f
C2510 a_244_55214# a_244_54862# 0.0109f
C2511 a_n908_55214# xaa0.xa2a.MN0.G 7.12e-19
C2512 xaa6.xe.XA7.MN1.G a_33652_54510# 7.1e-20
C2513 xaa6.xe.XA7.MP1.G a_32284_54510# 0.0969f
C2514 xaa0.xa1.MN0.G a_244_54158# 2.33e-19
C2515 xaa1.xa4.M0.D m3_37668_95644# 0.074f
C2516 xaa3.xa7.MN0.D a_4692_63422# 0.0972f
C2517 a_n908_63622# a_n908_63270# 0.0109f
C2518 xaa1.xa3.D xaa1.xa2.M6.D 0.00403f
C2519 a_4692_63774# xaa3.xa1b.MN0.D 7.59e-19
C2520 PWRUP_1V8 xaa6.xc.XA7.MN1.G 0.671f
C2521 AVDD xaa6.xc.XA7.MN0.D 0.485f
C2522 m2_4468_100124# m3_37748_100444# 0.0138f
C2523 xaa6.xd.XA1.MN0.G xaa6.xd.XA4.MN0.D 0.00303f
C2524 a_n908_55566# a_n908_55214# 0.0109f
C2525 xaa1.xa4.M0.D li_4468_103804# 23f
C2526 PWRUP_1V8 a_36172_54158# 0.00514f
C2527 a_26092_57326# xaa6.xc.XA5.MN0.G 6.98e-20
C2528 a_244_55566# xaa0.xa3.MP0.D 0.00176f
C2529 xaa0.xa1.MN0.G a_244_55214# 0.00329f
C2530 AVDD xaa0.xa1.MP1.D 0.191f
C2531 xaa3.xa3a.MN0.D li_6204_57236# 1.13e-19
C2532 a_4692_60078# li_4980_58996# 4.95e-20
C2533 CK m1_37504_57930# 0.0386f
C2534 a_29764_54862# a_31132_54862# 8.89e-19
C2535 xaa6.xg.XA4.MN0.G a_36172_54862# 0.0658f
C2536 a_37324_55214# a_37324_54862# 0.0109f
C2537 xaa1.xa4.M0.D m3_37748_112924# 0.111f
C2538 a_36172_52750# a_37324_52750# 0.00133f
C2539 xaa1.xa4.M0.D a_2948_74698# 0.383f
C2540 li_4468_70364# li_4468_70204# 7.91f
C2541 li_4468_90524# m1_4468_90524# 23f
C2542 PWRUP_1V8 xaa0.xa2a.MN0.D 0.579f
C2543 xaa5.xb1.MN1.D a_28612_61102# 0.0441f
C2544 AVDD a_27244_61102# 0.363f
C2545 m2_4468_113564# m3_37668_113884# 0.0138f
C2546 a_n76_76898# a_788_76898# 0.107f
C2547 xaa6.xg.XA7.MN1.G a_36172_56974# 0.00922f
C2548 IBPSR_1U xaa4.xa1.M6.D 0.026f
C2549 xaa6.xd.XA1.MN0.G xaa6.xd.XA6.MN0.D 0.00286f
C2550 xaa6.xe.XA7.MN1.G a_31132_56622# 0.0111f
C2551 xaa0.xa3.MN1.G a_244_56270# 0.00401f
C2552 a_n908_56622# a_n908_56270# 0.0109f
C2553 AVDD a_244_53806# 0.384f
C2554 xaa6.xf.XA6.MN0.G a_34804_54862# 0.0674f
C2555 xaa0.xa2a.MN0.G a_244_54510# 0.0896f
C2556 a_28612_55566# xaa6.xd.XA4.MP0.D 0.00176f
C2557 xaa1.xa4.M0.D m2_4468_116444# 71.5f
C2558 xaa6.xf.XA7.MN1.G a_33652_53102# 0.00893f
C2559 xaa6.xf.XA7.MP1.G a_34804_53102# 1.1e-19
C2560 xaa1.xa4.M0.D m3_4628_79164# 0.0276f
C2561 IBPSR_1U PWRUP_1V8 2.41f
C2562 xaa5.xb2_3.MN0.D CK 7.29e-20
C2563 a_27244_62862# a_28612_62862# 8.89e-19
C2564 AVDD xaa5.xb1.MN1.G 0.635f
C2565 m1_4468_90524# m2_4468_90524# 12.9f
C2566 xaa0.xa2a.MN0.D xaa0.xa5.MP1.D 1.28e-19
C2567 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN1.G 0.195f
C2568 a_36172_58030# xaa6.xg.XA7.MN1.G 8.24e-19
C2569 a_32284_57678# a_33652_57678# 8.89e-19
C2570 a_26092_57678# xaa6.xc.XA7.MN1.G 0.0736f
C2571 AVDD a_4692_55854# 0.00171f
C2572 m2_4468_86684# m3_37748_87004# 0.0138f
C2573 xaa6.xg.XA7.MN1.D a_37324_54158# 0.0747f
C2574 PWRUP_1V8 a_4308_51918# 4.07e-19
C2575 xaa6.xg.XA7.MP1.G xaa6.xg.XA3.MN0.D 0.0472f
C2576 xaa6.xg.XA7.MN1.G xaa6.xg.XA3.MP0.D 0.00242f
C2577 xaa6.xe.XA6.MN0.G a_32284_55918# 0.113f
C2578 xaa6.xe.XA7.MN1.G a_32284_54510# 0.0057f
C2579 xaa6.xe.XA7.MP1.G a_31132_54510# 0.0278f
C2580 xaa0.xa1.MN0.G a_n908_54158# 0.00564f
C2581 a_26092_55918# a_27244_55918# 0.00133f
C2582 a_28612_54158# a_29764_54158# 0.00133f
C2583 a_10092_54510# xaa4.xa1.M2.D 8.62e-20
C2584 xaa1.xa4.M0.D m3_4788_96444# 0.0138f
C2585 li_4468_104764# li_4468_103964# 39.3f
C2586 a_29764_64270# a_29764_63918# 0.0109f
C2587 xaa5.xb3.MP1.D a_28612_63566# 2.11e-19
C2588 AVDD xaa6.xc.XA7.MP1.G 2.06f
C2589 m2_4468_100124# m3_37668_100444# 0.0138f
C2590 xaa6.xd.XA1.MN0.G xaa6.xd.XA4.MP0.D 4.75e-19
C2591 xaa6.xd.XA7.MN1.D xaa6.xd.XA4.MN0.D 0.026f
C2592 PWRUP_1V8 a_34804_54158# 0.00514f
C2593 xaa0.xa1.MN0.G a_n908_55214# 0.0839f
C2594 a_29764_56622# xaa6.xd.XA6.MN0.D 0.00176f
C2595 xaa6.xd.XA7.MN1.G a_29764_55566# 7.66e-19
C2596 AVDD a_37324_54158# 0.386f
C2597 xaa3.xa3a.MN0.D li_6132_57236# 5.63e-20
C2598 a_4692_60078# li_4836_58996# 9.91e-20
C2599 a_5844_60078# li_6204_59524# 5.99e-19
C2600 xaa1.xa4.M0.D m3_37668_112924# 0.074f
C2601 a_2084_74698# a_2948_74698# 0.00813f
C2602 xaa1.xa1.M7.D xaa0.xa2a.MN0.D 0.00551f
C2603 PWRUP_1V8 xaa1.xa1.M5.D 5.67e-19
C2604 a_27244_61454# xaa5.xa3.xc1a.D 0.00176f
C2605 AVDD a_26092_61102# 0.00159f
C2606 xaa6.xd.XA7.MN1.D xaa6.xd.XA6.MN0.D 0.0989f
C2607 xaa6.xd.XA1.MN0.G xaa6.xd.XA6.MP0.D 4.47e-19
C2608 xaa0.xa3.MN1.G a_n908_56270# 0.0311f
C2609 a_244_56622# xaa0.xa5.MN0.D 0.0658f
C2610 a_n908_56622# xaa0.xa5.MN2.D 0.00176f
C2611 a_34804_57326# xaa6.xf.XA7.MN2.D 0.00176f
C2612 a_28612_57326# a_28612_56974# 0.0109f
C2613 IBPSR_1U a_11712_54334# 6.4e-19
C2614 AVDD a_n908_53806# 0.00159f
C2615 m2_4468_73244# m3_37748_73564# 0.0138f
C2616 xaa6.xf.XA5.MN0.G xaa6.xf.XA4.MN0.D 0.126f
C2617 xaa6.xf.XA6.MN0.G a_33652_54862# 0.0709f
C2618 xaa0.xa2a.MN0.G a_n908_54510# 0.112f
C2619 a_244_54862# a_244_54510# 0.0109f
C2620 xaa1.xa4.M0.D m2_4468_117404# 71.5f
C2621 a_10092_55566# a_10092_55038# 0.00702f
C2622 a_34804_53806# a_34804_53454# 0.0109f
C2623 xaa1.xa4.M0.D m3_37748_79324# 0.111f
C2624 li_4468_87644# li_4468_87484# 7.91f
C2625 li_4468_113564# m1_4468_113564# 23f
C2626 xaa5.xa3.xb2_0.G a_27244_61806# 7.73e-19
C2627 IBPSR_1U xaa1.xa1.M7.D 0.026f
C2628 xaa5.xb1.MN1.G xaa5.xb1.MN1.D 0.209f
C2629 a_29764_63214# CK 3.97e-20
C2630 xaa5.xb2_3.MN0.D a_29764_62862# 0.126f
C2631 AVDD xaa3.xa1b.MN0.D 1.4f
C2632 xaa6.xd.XA7.MN1.D xaa6.xe.XA7.MN1.G 7.59e-20
C2633 xaa6.xe.XA7.MN1.D xaa6.xd.XA7.MN1.G 7.59e-20
C2634 AVDD a_5844_56206# 0.348f
C2635 m2_4468_86684# m3_37668_87004# 0.0138f
C2636 xaa6.xg.XA7.MN1.D a_36172_54158# 0.066f
C2637 xaa6.xf.XA1.MN0.G a_37324_54158# 1.11e-19
C2638 xaa6.xg.XA7.MP1.G xaa6.xg.XA3.MN1.G 0.352f
C2639 xaa6.xe.XA6.MN0.G a_31132_55918# 0.0873f
C2640 a_36172_56270# a_36172_55918# 0.0109f
C2641 xaa0.xa3.MP0.D a_244_54862# 0.00176f
C2642 a_n908_55214# a_n908_54862# 0.0109f
C2643 xaa6.xe.XA7.MN1.G a_31132_54510# 0.082f
C2644 a_26092_56270# xaa6.xc.XA5.MN0.G 0.00131f
C2645 a_37324_54510# a_37324_54158# 0.0109f
C2646 xaa1.xa4.M0.D m3_4628_96444# 0.0276f
C2647 xaa3.xa7.MN0.D xaa3.xa8.MP0.D 0.01f
C2648 xaa0.xa6.MN0.D xaa1.xa2.M8.D 0.0176f
C2649 xaa5.xb3.MP1.D xaa5.xa3.xb2_0.G 6.83e-19
C2650 a_5844_63774# a_5844_63422# 0.0109f
C2651 li_4468_69404# m1_4468_69404# 23f
C2652 xaa0.xa6.MN0.D xaa0.xa3.MP0.D 3.47e-20
C2653 xaa4.xa4.M0.D a_11712_59086# 0.154f
C2654 a_n908_59750# a_640_59750# 6.96e-19
C2655 AVDD xaa6.xc.XA7.MN1.G 3.53f
C2656 xaa6.xf.XA7.MN1.G xaa6.xf.XA5.MN0.G 0.0911f
C2657 xaa6.xc.XA1.MN0.G xaa6.xd.XA4.MN0.D 3.2e-19
C2658 xaa6.xd.XA7.MN1.D xaa6.xd.XA4.MP0.D 0.00426f
C2659 a_n908_55566# a_244_55566# 0.00133f
C2660 xaa1.xa4.M0.D li_4468_104764# 23f
C2661 xaa0.xa1.MN0.G xaa0.xa3.MP0.D 0.0624f
C2662 xaa6.xd.XA7.MP1.G a_29764_55566# 0.0964f
C2663 xaa6.xd.XA7.MN1.G a_28612_55566# 0.0769f
C2664 AVDD a_36172_54158# 0.00156f
C2665 xaa3.xa3a.MN0.D li_4980_58996# 0.0249f
C2666 a_5844_60078# li_6132_59524# 2e-19
C2667 a_28612_54862# a_29764_54862# 0.00133f
C2668 a_36172_55214# a_36172_54862# 0.0109f
C2669 a_2948_70022# m2_4468_69404# 3.37e-19
C2670 xaa1.xa4.M0.D m3_4788_113724# 0.0138f
C2671 a_34804_52750# a_36172_52750# 8.89e-19
C2672 li_4468_71164# li_4468_70364# 39.3f
C2673 PWRUP_1V8 xaa5.xb1.MN0.D 0.0111f
C2674 xaa1.xa1.M8.D xaa0.xa2a.MN0.D 0.0984f
C2675 CK a_29764_60750# 1.02e-20
C2676 a_n508_74698# a_356_74698# 0.071f
C2677 AVDD xaa0.xa2a.MN0.D 1.72f
C2678 xaa6.xc.XA1.MN0.G xaa6.xd.XA6.MN0.D 3e-19
C2679 xaa6.xd.XA7.MN1.D xaa6.xd.XA6.MP0.D 0.0532f
C2680 xaa6.xd.XA7.MN0.D a_29764_56622# 1.28e-19
C2681 a_n908_56622# xaa0.xa5.MN0.D 0.0677f
C2682 xaa0.xa3.MN1.G xaa0.xa5.MN2.D 0.152f
C2683 xaa6.xf.XA7.MN0.D a_34804_56974# 0.00297f
C2684 IBPSR_1U xaa4.xa1.M7.D 0.026f
C2685 AVDD xaa0.xa1.MN2.D 0.00193f
C2686 m2_4468_73244# m3_37668_73564# 0.0138f
C2687 xaa6.xf.XA5.MN0.G xaa6.xf.XA4.MP0.D 0.0618f
C2688 a_27244_55566# xaa6.xc.XA4.MP0.D 0.00176f
C2689 xaa6.xc.XA7.MN1.G a_27244_52750# 0.00154f
C2690 xaa1.xa4.M0.D m3_37668_79324# 0.074f
C2691 xaa4.xa2.M0.G a_29764_61806# 3.48e-19
C2692 IBPSR_1U xaa1.xa1.M8.D 0.0482f
C2693 xaa5.xa3.xb2_0.G a_26092_61806# 0.175f
C2694 xaa1.xa3.D xaa1.xb2.M0.D 0.00297f
C2695 xaa0.xa6.MN0.D xaa1.xa1.M6.D 6.39e-19
C2696 a_29764_63214# a_29764_62862# 0.0109f
C2697 xaa5.xb2_3.MN0.D a_28612_62862# 0.0878f
C2698 a_26092_62862# a_27244_62862# 0.00133f
C2699 AVDD IBPSR_1U 1.84f
C2700 m1_4468_91484# m2_4468_91484# 12.9f
C2701 xaa6.xd.XA1.MN0.G xaa6.xd.XA7.MN1.G 0.224f
C2702 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MN0.D 0.336f
C2703 a_31132_57678# a_32284_57678# 0.00133f
C2704 AVDD a_4692_56206# 0.00171f
C2705 xaa0.xa5.MN2.G a_244_52750# 2.36e-19
C2706 xaa6.xf.XA1.MN0.G a_36172_54158# 0.00207f
C2707 xaa6.xg.XA7.MN1.G xaa6.xg.XA3.MN1.G 0.129f
C2708 xaa0.xa1.MN0.G a_n908_54510# 0.0046f
C2709 xaa4.xa4.M0.D xaa4.xa1.M1.D 4.85e-19
C2710 a_27244_54158# a_28612_54158# 8.89e-19
C2711 xaa1.xa4.M0.D m3_37748_96604# 0.111f
C2712 li_4468_104924# li_4468_104764# 7.91f
C2713 a_n908_63622# xaa1.xa2.M8.D 0.00224f
C2714 a_28612_64270# a_28612_63918# 0.0109f
C2715 a_29764_64270# xaa4.xa2.M0.G 3.48e-19
C2716 xaa1.xa3.D xaa1.xa2.M7.D 0.00622f
C2717 xaa0.xa6.MN0.D a_244_55566# 5.27e-19
C2718 PWRUP_1V8 a_36172_57678# 0.0042f
C2719 a_11712_60670# a_11712_59086# 0.00223f
C2720 xaa3.xa3a.MN0.D a_5844_57790# 7.03e-19
C2721 AVDD a_11712_57502# 0.424f
C2722 xaa6.xf.XA7.MP1.G xaa6.xf.XA5.MN0.G 0.397f
C2723 xaa6.xc.XA1.MN0.G xaa6.xd.XA4.MP0.D 0.00287f
C2724 xaa0.xa1.MN0.G a_244_55566# 0.0889f
C2725 a_28612_56622# xaa6.xd.XA6.MP0.D 0.00176f
C2726 xaa6.xd.XA7.MP1.G a_28612_55566# 0.0292f
C2727 xaa6.xd.XA7.MN1.G a_27244_55566# 7.1e-20
C2728 xaa6.xf.XA7.MN1.G xaa6.xe.XA5.MN0.G 1.74e-19
C2729 AVDD a_34804_54158# 0.00156f
C2730 a_2948_70022# m2_4468_70364# 0.00238f
C2731 xaa1.xa4.M0.D m3_4628_113724# 0.0276f
C2732 xaa3.xa3a.MN0.D li_4836_58996# 0.0139f
C2733 a_2084_74698# xaa1.xa4.M0.D 0.0492f
C2734 li_4468_91484# m1_4468_91484# 23f
C2735 xaa1.xa1.M8.D xaa1.xa1.M5.D 0.00345f
C2736 xaa5.xa3.xb2_0.D a_27244_60750# 0.071f
C2737 a_28612_61454# a_29764_61454# 0.00133f
C2738 xbb0.xa1.XA1.N a_788_76898# 0.00114f
C2739 xaa6.xc.XA1.MN0.G xaa6.xd.XA6.MP0.D 0.00276f
C2740 xaa6.xd.XA7.MN0.D a_28612_56622# 0.0217f
C2741 xaa6.xd.XA7.MN1.G a_29764_56622# 0.0111f
C2742 a_n908_56622# a_244_56622# 0.00133f
C2743 xaa0.xa3.MN1.G xaa0.xa5.MN0.D 0.446f
C2744 a_27244_57326# a_27244_56974# 0.0109f
C2745 xaa6.xf.XA7.MN1.G a_34804_56974# 0.00922f
C2746 xaa6.xf.XA7.MN0.D a_33652_56974# 0.016f
C2747 AVDD xaa0.xa1.MN0.D 0.702f
C2748 xaa6.xe.XA6.MN0.G a_32284_54862# 0.0725f
C2749 a_244_54862# xaa0.xa2a.MN0.G 0.0658f
C2750 a_n908_54862# a_n908_54510# 0.0109f
C2751 xaa6.xc.XA7.MN1.G a_26092_52750# 2.64e-19
C2752 a_4692_62366# li_4980_61284# 4.95e-20
C2753 xaa3.xa5a.MN0.D li_6204_59524# 1.13e-19
C2754 xaa6.xc.XA1.MN0.D a_26092_53454# 0.0492f
C2755 a_33652_53806# a_33652_53454# 0.0109f
C2756 xaa1.xa4.M0.D m3_4788_80124# 0.0138f
C2757 li_4468_88444# li_4468_87644# 39.3f
C2758 xaa4.xa2.M0.G a_28612_61806# 0.0362f
C2759 a_27244_63214# CK 0.0021f
C2760 AVDD a_n908_63270# 7.8e-20
C2761 m1_37504_57930# m1_37504_55818# 0.00656f
C2762 xaa6.xd.XA1.MN0.G xaa6.xd.XA7.MP1.G 0.0184f
C2763 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN0.D 0.129f
C2764 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MN1.G 0.467f
C2765 xaa6.xg.XA7.MN1.D a_37324_57678# 0.0893f
C2766 a_34804_58030# xaa6.xf.XA7.MN1.G 0.00227f
C2767 AVDD xaa0.xa1.MN2.S 1.24f
C2768 xaa6.xf.XA1.MN0.G a_34804_54158# 0.00268f
C2769 xaa0.xa5.MN2.G a_n908_52750# 2.76e-19
C2770 xaa6.xd.XA6.MN0.G a_29764_55918# 0.0889f
C2771 a_34804_56270# a_34804_55918# 0.0109f
C2772 xaa0.xa1.MN0.G xaa0.xa2a.MN0.G 0.0982f
C2773 a_36172_54510# a_36172_54158# 0.0109f
C2774 xaa1.xa4.M0.D m3_37668_96604# 0.074f
C2775 a_28612_64270# xaa4.xa2.M0.G 0.0138f
C2776 a_29764_64270# xaa5.xa3.xb1_0.G 0.0701f
C2777 xaa1.xa4.M0.G xaa3.xa1b.MN0.D 0.0387f
C2778 xaa5.xb3.MP1.D a_28612_63918# 6.57e-19
C2779 a_4692_63774# a_4692_63422# 0.0109f
C2780 li_4468_70204# m1_4468_70204# 23f
C2781 CK a_37324_57326# 5.74e-19
C2782 PWRUP_1V8 a_34804_57678# 0.00444f
C2783 xaa3.xa3a.MN0.D a_4692_57790# 1.15e-19
C2784 xaa0.xa6.MN0.D a_n908_55566# 8.92e-20
C2785 AVDD a_37324_57678# 0.383f
C2786 xaa6.xc.XA1.MN0.G xaa6.xc.XA4.MP0.D 0.00303f
C2787 xaa1.xa4.M0.D li_4468_105724# 23f
C2788 PWRUP_1V8 a_31132_54158# 0.00514f
C2789 xaa0.xa1.MN0.G a_n908_55566# 0.0794f
C2790 a_244_55918# a_244_55566# 0.0109f
C2791 AVDD a_33652_54158# 0.387f
C2792 a_27244_54862# a_28612_54862# 8.89e-19
C2793 a_34804_55214# a_34804_54862# 0.0109f
C2794 a_2948_70022# m2_4468_71324# 0.00238f
C2795 xaa1.xa3.D m2_4468_69404# 59.5f
C2796 xaa1.xa4.M0.D m3_37748_113884# 0.111f
C2797 xaa3.xa3a.MN0.D li_6204_59524# 0.118f
C2798 a_33652_52750# a_34804_52750# 0.00133f
C2799 xaa6.xg.XA6.MN0.G m1_37504_55818# 0.0501f
C2800 a_1652_76898# a_2948_74698# 0.00121f
C2801 li_4468_71324# li_4468_71164# 7.91f
C2802 PWRUP_1V8 a_640_61158# 0.0744f
C2803 xaa5.xa3.xb2_0.D a_26092_60750# 3.3e-20
C2804 AVDD xaa5.xb1.MN0.D 4.89e-20
C2805 a_n940_74698# a_788_76898# 2.35e-20
C2806 xbb0.xa1.XA1.N a_356_74698# 0.00388f
C2807 m2_4468_114524# m3_37748_114844# 0.0138f
C2808 xaa6.xc.XA1.MN0.G xaa6.xc.XA6.MP0.D 0.00286f
C2809 xaa6.xd.XA7.MN1.G a_28612_56622# 0.0785f
C2810 xaa6.xd.XA7.MP1.G a_29764_56622# 0.0676f
C2811 xaa0.xa3.MN1.G a_244_56622# 0.0896f
C2812 xaa6.xf.XA7.MP1.G a_34804_56974# 2.35e-19
C2813 xaa6.xf.XA7.MN1.G a_33652_56974# 0.0035f
C2814 xaa4.xa4.M0.D a_11712_55918# 0.0877f
C2815 AVDD a_244_54158# 0.388f
C2816 a_n908_54862# xaa0.xa2a.MN0.G 0.0731f
C2817 a_26092_55566# xaa6.xc.XA4.MN0.D 0.00176f
C2818 xaa6.xe.XA5.MN0.G xaa6.xe.XA4.MP0.D 0.0618f
C2819 a_4692_62366# li_4836_61284# 9.91e-20
C2820 a_5844_62366# li_6204_61812# 5.99e-19
C2821 xaa3.xa5a.MN0.D li_6132_59524# 5.63e-20
C2822 xaa6.xe.XA6.MN0.G a_31132_54862# 0.0658f
C2823 xaa1.xa4.M0.D m3_4628_80124# 0.0276f
C2824 li_4468_114524# m1_4468_114524# 23f
C2825 xaa4.xa2.M0.G a_27244_61806# 5.56e-19
C2826 xaa5.xa3.xb2_0.G xaa5.xb2_0.MN0.D 0.00104f
C2827 xaa5.xb1.MN1.G a_29764_61806# 0.00688f
C2828 a_26092_63214# CK 0.00969f
C2829 a_28612_63214# a_28612_62862# 0.0109f
C2830 AVDD a_5844_63422# 0.364f
C2831 m1_4468_92444# m2_4468_92444# 12.9f
C2832 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN1.G 0.201f
C2833 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MP1.G 0.313f
C2834 a_29764_57678# a_31132_57678# 8.89e-19
C2835 xaa6.xg.XA7.MN1.D a_36172_57678# 0.132f
C2836 xaa6.xf.XA1.MN0.G a_37324_57678# 0.00235f
C2837 a_33652_58030# xaa6.xf.XA7.MN1.G 1.55e-20
C2838 AVDD a_244_55214# 0.364f
C2839 xaa6.xd.XA7.MN1.G a_29764_54510# 0.0835f
C2840 xaa6.xf.XA1.MN0.G a_33652_54158# 1.35e-19
C2841 xaa6.xf.XA7.MN1.D a_34804_54158# 0.0676f
C2842 xaa6.xd.XA6.MN0.G a_28612_55918# 0.111f
C2843 xaa0.xa1.MN0.G a_244_54862# 3.61e-19
C2844 xaa6.xf.XA7.MN1.G xaa6.xg.XA3.MN1.G 0.00435f
C2845 a_26092_54158# a_27244_54158# 0.00133f
C2846 xaa1.xa4.M0.D m3_4788_97404# 0.0138f
C2847 li_4468_105724# li_4468_104924# 39.3f
C2848 xaa5.xb3.MP1.D xaa4.xa2.M0.G 0.0548f
C2849 a_28612_64270# xaa5.xa3.xb1_0.G 0.07f
C2850 a_29764_64270# xaa5.xb1.MN1.G 0.0309f
C2851 xaa1.xa4.M0.G IBPSR_1U 4.6e-19
C2852 a_5844_63774# xaa3.xa8.MP0.D 0.00176f
C2853 xaa3.xa3a.MN0.D xaa3.xa1capd.B 0.00369f
C2854 xaa0.xa6.MN0.D xaa0.xa1.MN0.G 0.00263f
C2855 AVDD a_36172_57678# 0.00163f
C2856 m2_4468_101084# m3_37748_101404# 0.0138f
C2857 xaa6.xc.XA1.MN0.G xaa6.xc.XA4.MN0.D 4.75e-19
C2858 PWRUP_1V8 a_29764_54158# 0.00514f
C2859 xaa6.xc.XA7.MN1.D xaa6.xc.XA4.MP0.D 0.00426f
C2860 a_27244_56622# xaa6.xc.XA6.MP0.D 0.00176f
C2861 AVDD a_32284_54158# 0.387f
C2862 a_2948_70022# m2_4468_72284# 0.00125f
C2863 xaa1.xa3.D m2_4468_70364# 71.5f
C2864 xaa1.xa4.M0.D m3_37668_113884# 0.074f
C2865 xaa3.xa3a.MN0.D li_6132_59524# 0.0319f
C2866 a_1220_74698# a_2948_74698# 9.03e-19
C2867 PWRUP_1V8 xaa1.xa1.M6.D 0.00538f
C2868 xaa5.xb1.MN1.D xaa5.xb1.MN0.D 0.106f
C2869 a_27244_61454# a_28612_61454# 8.89e-19
C2870 a_n908_61510# xaa0.xa2a.MN0.D 4.86e-19
C2871 AVDD xaa5.xa3.xc1a.D 0.153f
C2872 a_n940_74698# a_356_74698# 9.03e-19
C2873 m2_4468_114524# m3_37668_114844# 0.0138f
C2874 xaa6.xc.XA1.MN0.G xaa6.xc.XA6.MN0.D 4.47e-19
C2875 xaa6.xd.XA7.MP1.G a_28612_56622# 0.029f
C2876 xaa0.xa3.MN1.G a_n908_56622# 0.0885f
C2877 a_244_56974# a_244_56622# 0.0109f
C2878 a_31132_57326# xaa6.xe.XA7.MN2.D 0.00176f
C2879 a_26092_57326# a_26092_56974# 0.0109f
C2880 a_n908_56974# xaa0.xa5.MN0.D 1.21e-19
C2881 xaa6.xf.XA7.MP1.G a_33652_56974# 0.0291f
C2882 xaa6.xc.XA7.MN1.D xaa6.xc.XA6.MP0.D 0.0532f
C2883 AVDD a_n908_54158# 0.00171f
C2884 xaa6.xe.XA7.MP1.G a_31132_53102# 1.1e-19
C2885 xaa6.xe.XA7.MN1.G a_32284_53102# 0.00893f
C2886 a_n908_54862# a_244_54862# 0.00133f
C2887 xaa6.xe.XA5.MN0.G xaa6.xe.XA4.MN0.D 0.126f
C2888 a_5844_62366# li_6132_61812# 2e-19
C2889 xaa3.xa5a.MN0.D li_4980_61284# 0.0249f
C2890 a_32284_53806# a_32284_53454# 0.0109f
C2891 xbb1.xa3.M6.D xbb1.xa3.M5.D 0.0488f
C2892 xaa1.xa4.M0.D m3_37748_80284# 0.111f
C2893 li_4468_88604# li_4468_88444# 7.91f
C2894 IBPSR_1U a_n908_61510# 0.156f
C2895 xaa5.xa3.xb2_0.G xaa5.xa3.xc2a.D 0.00186f
C2896 xaa5.xb1.MN1.G a_28612_61806# 9.6e-19
C2897 AVDD a_4692_63422# 0.00159f
C2898 xaa6.xc.XA7.MN1.D xaa6.xd.XA7.MN1.G 1.74e-19
C2899 xaa4.xa2.M0.G xaa4.xa1.M8.D 0.0709f
C2900 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MP1.G 0.216f
C2901 AVDD a_n908_55214# 0.00159f
C2902 xaa6.xf.XA1.MN0.G a_36172_57678# 0.00674f
C2903 a_33652_58030# xaa6.xf.XA7.MP1.G 3.8e-19
C2904 m2_4468_87644# m3_37748_87964# 0.0138f
C2905 xaa6.xd.XA7.MN1.G a_28612_54510# 0.0057f
C2906 xaa6.xd.XA7.MP1.G a_29764_54510# 0.0278f
C2907 xaa6.xe.XA1.MN0.G a_34804_54158# 1.11e-19
C2908 xaa6.xf.XA7.MN1.D a_33652_54158# 0.0731f
C2909 xaa0.xa5.MN2.G a_n908_53102# 4.05e-20
C2910 a_33652_56270# a_33652_55918# 0.0109f
C2911 xaa0.xa1.MN0.G a_n908_54862# 0.0106f
C2912 xaa6.xf.XA7.MN1.G xaa6.xf.XA3.MN0.D 0.0288f
C2913 a_34804_54510# a_34804_54158# 0.0109f
C2914 xaa1.xa4.M0.D m3_4628_97404# 0.0276f
C2915 xaa6.xg.XA4.MN0.G m1_37504_55818# 0.0493f
C2916 a_28612_64270# xaa5.xb1.MN1.G 0.0215f
C2917 xaa1.xa4.M0.G a_n908_63270# 2.92e-19
C2918 xaa5.xb3.MP1.D xaa5.xa3.xb1_0.G 0.0258f
C2919 a_29764_64622# xaa4.xa2.M0.G 0.00113f
C2920 a_5844_63774# xaa3.xa7.MN0.D 0.0658f
C2921 a_n908_63622# xaa0.xa6.MN0.D 0.0725f
C2922 li_4468_70364# m1_4468_70364# 23f
C2923 a_11712_60670# xaa4.xa4.M0.D 0.0676f
C2924 xaa3.xa3a.MN0.D a_5844_58142# 0.00414f
C2925 a_5844_60078# a_5844_58494# 0.00744f
C2926 xaa0.xa6.MN0.D a_244_55918# 8.96e-19
C2927 AVDD a_34804_57678# 0.00163f
C2928 m2_4468_101084# m3_37668_101404# 0.0138f
C2929 xaa1.xa4.M0.D li_4468_106684# 23f
C2930 IBPSR_1U a_10092_52750# 0.0705f
C2931 xaa3.xa1b.MN0.D xbb1.xa3.M3.D 1.38e-19
C2932 a_n908_55918# a_n908_55566# 0.0109f
C2933 xaa6.xc.XA7.MN1.G a_28612_55566# 7.1e-20
C2934 xaa6.xc.XA7.MP1.G a_27244_55566# 0.0292f
C2935 xaa6.xe.XA7.MP1.G xaa6.xe.XA5.MN0.G 0.397f
C2936 xaa6.xc.XA7.MN1.D xaa6.xc.XA4.MN0.D 0.026f
C2937 xaa0.xa5.MP1.D a_244_55566# 0.00176f
C2938 xaa6.xe.XA7.MN1.G xaa6.xf.XA5.MN0.G 1.74e-19
C2939 a_244_55918# xaa0.xa1.MN0.G 0.0661f
C2940 AVDD a_31132_54158# 0.00156f
C2941 a_26092_54862# a_27244_54862# 0.00133f
C2942 a_33652_55214# a_33652_54862# 0.0109f
C2943 xaa1.xa3.D m2_4468_71324# 71.5f
C2944 xaa1.xa4.M0.D m3_4788_114684# 0.0138f
C2945 a_32284_52750# a_33652_52750# 8.89e-19
C2946 a_1652_76898# xaa1.xa4.M0.D 0.163f
C2947 li_4468_72124# li_4468_71324# 39.3f
C2948 li_4468_92444# m1_4468_92444# 23f
C2949 PWRUP_1V8 a_29764_61454# 1.28e-19
C2950 xaa1.xa1.M7.D xaa1.xa1.M6.D 0.0488f
C2951 xaa1.xa1.M8.D a_640_61158# 0.0177f
C2952 a_n908_61510# xaa1.xa1.M5.D 2.99e-19
C2953 AVDD a_640_61158# 0.376f
C2954 AVDD a_244_54510# 0.388f
C2955 xaa6.xc.XA7.MN1.D xaa6.xc.XA6.MN0.D 0.0989f
C2956 xaa0.xa5.MN2.G xaa6.xc.XA6.MP0.D 4.24e-20
C2957 m2_4468_74204# m3_37748_74524# 0.0138f
C2958 xaa4.xa2.M0.D a_10092_55038# 0.00624f
C2959 xaa6.xe.XA7.MN1.G a_31132_53102# 7.44e-19
C2960 xaa6.xg.XA7.MN1.D a_37324_52750# 3.67e-21
C2961 xaa3.xa5a.MN0.D li_4836_61284# 0.0139f
C2962 xaa6.xg.XA7.MP1.G a_37324_53454# 1.07e-19
C2963 xaa6.xd.XA6.MN0.G a_29764_54862# 0.0674f
C2964 xaa1.xa4.M0.D m3_37668_80284# 0.074f
C2965 a_27244_63214# a_27244_62862# 0.0109f
C2966 a_29764_63214# xaa5.xb2_3.MN0.D 0.0682f
C2967 xaa1.xa3.D a_640_60806# 0.00485f
C2968 xaa5.xa3.xb1_0.G a_26092_61806# 0.00207f
C2969 m1_4468_93404# m2_4468_93404# 12.9f
C2970 xaa6.xc.XA1.MN0.G xaa6.xc.XA7.MN0.D 0.00664f
C2971 a_28612_57678# a_29764_57678# 0.00133f
C2972 xaa6.xf.XA1.MN0.G a_34804_57678# 0.00219f
C2973 AVDD xaa0.xa3.MP0.D 0.191f
C2974 m2_4468_87644# m3_37668_87964# 0.0138f
C2975 xaa6.xd.XA7.MP1.G a_28612_54510# 0.0953f
C2976 xaa6.xd.XA7.MN1.G a_27244_54510# 7.1e-20
C2977 xaa6.xe.XA1.MN0.G a_33652_54158# 0.00209f
C2978 xaa6.xf.XA6.MN0.G xaa6.xg.XA6.MN0.G 0.00217f
C2979 xaa6.xc.XA6.MN0.G a_27244_55918# 0.113f
C2980 xaa1.xa4.M0.D li_4468_73084# 23f
C2981 PWRUP_1V8 a_34804_52750# 4.95e-20
C2982 xaa6.xf.XA7.MP1.G xaa6.xf.XA3.MN0.D 0.0472f
C2983 xaa6.xf.XA7.MN1.G xaa6.xf.XA3.MP0.D 0.00252f
C2984 AVDD a_37324_52750# 0.448f
C2985 xaa1.xa4.M0.D m3_37748_97564# 0.111f
C2986 a_37324_55214# m1_37504_55818# 0.0137f
C2987 li_4468_105884# li_4468_105724# 7.91f
C2988 a_28612_64622# xaa4.xa2.M0.G 0.0123f
C2989 xaa1.xa4.M0.G a_5844_63422# 0.00276f
C2990 xaa5.xb3.MP1.D xaa5.xb1.MN1.G 0.0424f
C2991 a_29764_64622# xaa5.xa3.xb1_0.G 1.75e-19
C2992 a_4692_63774# xaa3.xa7.MN0.D 0.0711f
C2993 PWRUP_1V8 a_31132_57678# 0.0042f
C2994 xaa3.xa3a.MN0.D a_4692_58142# 0.00348f
C2995 xaa0.xa6.MN0.D a_n908_55918# 1.52e-19
C2996 AVDD a_33652_57678# 0.384f
C2997 AVDD a_29764_54158# 0.00156f
C2998 IBPSR_1U xbb1.xa3.M3.D 0.0497f
C2999 xaa6.xc.XA7.MN1.G a_27244_55566# 0.0754f
C3000 xaa6.xc.XA7.MP1.G a_26092_55566# 0.098f
C3001 xaa6.xe.XA7.MN1.G xaa6.xe.XA5.MN0.G 0.0911f
C3002 CK a_36172_53806# 1.32e-19
C3003 a_26092_56622# xaa6.xc.XA6.MN0.D 0.00176f
C3004 a_n908_55918# xaa0.xa1.MN0.G 0.065f
C3005 xaa1.xa3.D m2_4468_72284# 12f
C3006 xaa1.xa4.M0.D m3_4628_114684# 0.0276f
C3007 xbb1.xa3.M3.D a_4308_51918# 1.81e-19
C3008 a_1220_74698# xaa1.xa4.M0.D 0.00282f
C3009 xaa1.xa1.M8.D xaa1.xa1.M6.D 0.00611f
C3010 a_26092_61454# a_27244_61454# 0.00133f
C3011 xaa4.xa2.M0.G xaa0.xa5.MN2.G 0.0248f
C3012 xbb0.xa1.XA1.N a_n76_76898# 0.119f
C3013 xaa6.xc.XA7.MN0.D a_27244_56622# 0.0217f
C3014 a_244_56974# xaa0.xa3.MN1.G 0.0658f
C3015 a_n908_56974# a_n908_56622# 0.0109f
C3016 a_29764_57326# xaa6.xd.XA7.MN2.D 0.00176f
C3017 xaa6.xg.XA7.MN0.D xaa6.xg.XA7.MN2.D 0.0618f
C3018 xaa6.xe.XA7.MN0.D a_32284_56974# 0.016f
C3019 AVDD a_n908_54510# 0.00171f
C3020 m2_4468_74204# m3_37668_74524# 0.0138f
C3021 xaa6.xg.XA7.MN1.D a_36172_52750# 6.12e-22
C3022 xaa6.xd.XA5.MN0.G xaa6.xd.XA4.MN0.D 0.126f
C3023 xaa3.xa5a.MN0.D li_6204_61812# 0.118f
C3024 xaa6.xg.XA7.MN1.G a_37324_53454# 0.0204f
C3025 xaa6.xg.XA7.MP1.G a_36172_53454# 2.78e-19
C3026 xaa6.xd.XA6.MN0.G a_28612_54862# 0.0709f
C3027 a_37324_57326# m1_37504_55818# 5e-20
C3028 a_31132_53806# a_31132_53454# 0.0109f
C3029 xaa4.xa1.M2.D xaa4.xa1.M1.D 0.0488f
C3030 xaa1.xa4.M0.D m3_4788_81084# 0.0138f
C3031 li_4468_115484# m1_4468_115484# 23f
C3032 li_4468_89404# li_4468_88604# 39.3f
C3033 xaa0.xa6.MN0.D PWRUP_1V8 0.181f
C3034 a_28612_63214# xaa5.xb2_3.MN0.D 0.0674f
C3035 xaa4.xa2.M0.G xaa5.xb2_0.MN0.D 0.174f
C3036 xaa5.xa3.xb2_0.G a_29764_62158# 1.11e-19
C3037 AVDD xaa3.xa8.MP0.D 0.191f
C3038 m1_4468_70204# m1_4468_69404# 56.4f
C3039 xaa0.xa5.MN2.G xaa6.xd.XA7.MP1.G 4.23e-19
C3040 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MN0.D 0.336f
C3041 xaa6.xc.XA1.MN0.G xaa6.xc.XA7.MP1.G 0.027f
C3042 PWRUP_1V8 xaa0.xa1.MN0.G 0.238f
C3043 xaa6.xd.XA7.MN1.D xaa6.xc.XA7.MN1.G 1.74e-19
C3044 xaa6.xf.XA7.MN1.D a_34804_57678# 0.134f
C3045 xaa6.xf.XA1.MN0.G a_33652_57678# 1.35e-19
C3046 AVDD a_244_55566# 0.383f
C3047 xaa6.xe.XA1.MN0.G a_32284_54158# 0.00329f
C3048 xaa0.xa5.MN2.G a_n908_53454# 4.05e-20
C3049 xaa6.xc.XA6.MN0.G a_26092_55918# 0.0873f
C3050 a_32284_56270# a_32284_55918# 0.0109f
C3051 AVDD a_36172_52750# 0.00535f
C3052 a_2948_74698# li_4468_74204# 1.18e-19
C3053 xaa6.xf.XA7.MP1.G xaa6.xf.XA3.MP0.D 0.0712f
C3054 xaa1.xa4.M0.D m3_37668_97564# 0.074f
C3055 a_33652_54510# a_33652_54158# 0.0109f
C3056 xaa1.xa4.M0.G a_4692_63422# 0.062f
C3057 a_29764_64622# xaa5.xb1.MN1.G 0.0012f
C3058 a_28612_64622# xaa5.xa3.xb1_0.G 0.00126f
C3059 xaa3.xa9.MN0.D xaa3.xa7.MN0.D 2.11e-19
C3060 li_4468_71164# m1_4468_71164# 23f
C3061 a_4692_60078# a_4692_58494# 0.00744f
C3062 xaa3.xa3a.MN0.D xaa3.xa2.MN0.D 0.175f
C3063 PWRUP_1V8 a_29764_57678# 0.00444f
C3064 xaa0.xa6.MN0.D xaa0.xa5.MP1.D 1.67e-19
C3065 AVDD a_32284_57678# 0.384f
C3066 xaa1.xa4.M0.D li_4468_107644# 23f
C3067 PWRUP_1V8 a_26092_54158# 0.00506f
C3068 xaa6.xc.XA7.MN1.G a_26092_55566# 7.66e-19
C3069 xaa0.xa5.MN2.G CK_REF 0.0353f
C3070 a_n908_55918# a_244_55918# 0.00133f
C3071 xaa0.xa5.MP1.D xaa0.xa1.MN0.G 0.0099f
C3072 AVDD a_28612_54158# 0.387f
C3073 a_32284_55214# a_32284_54862# 0.0109f
C3074 xaa1.xa4.M0.D m3_37748_114844# 0.111f
C3075 a_31132_52750# a_32284_52750# 0.00133f
C3076 a_1220_74698# a_2084_74698# 0.071f
C3077 li_4468_72284# li_4468_72124# 7.91f
C3078 a_640_61510# a_640_61158# 0.0109f
C3079 AVDD a_29764_61454# 0.00139f
C3080 a_n940_74698# a_n76_76898# 0.00121f
C3081 xbb0.xa1.XA1.N a_n508_74698# 0.207f
C3082 xaa6.xc.XA7.MN0.D a_26092_56622# 1.28e-19
C3083 xaa6.xe.XA7.MP1.G a_32284_56974# 0.0291f
C3084 xaa6.xg.XA7.MN0.D xaa6.xg.XA7.MN0.G 0.0903f
C3085 a_n908_56974# xaa0.xa3.MN1.G 0.0738f
C3086 xaa6.xc.XA7.MP1.G a_27244_56622# 0.029f
C3087 xaa6.xe.XA7.MN0.D a_31132_56974# 0.00297f
C3088 AVDD xaa0.xa2a.MN0.G 0.717f
C3089 xaa6.xd.XA5.MN0.G xaa6.xd.XA4.MP0.D 0.0618f
C3090 xaa3.xa5a.MN0.D li_6132_61812# 0.0319f
C3091 xaa6.xg.XA7.MN1.G a_36172_53454# 1.87e-19
C3092 xaa6.xf.XA6.MN0.G xaa6.xg.XA4.MN0.G 0.00217f
C3093 a_37324_57326# m1_37504_57930# 0.0134f
C3094 a_4308_53678# xbb1.xa3.M4.D 1.81e-19
C3095 xaa1.xa4.M0.D m3_4628_81084# 0.0276f
C3096 xaa0.xa6.MN0.D xaa1.xa1.M7.D 7.41e-19
C3097 a_26092_63214# a_26092_62862# 0.0109f
C3098 a_28612_63214# a_29764_63214# 0.00133f
C3099 xaa1.xa3.D xaa1.xb2.M7.D 0.076f
C3100 xaa5.xa3.xb2_0.G a_28612_62158# 5.27e-19
C3101 xaa4.xa2.M0.G xaa5.xa3.xc2a.D 1.46e-19
C3102 AVDD xaa3.xa7.MN0.D 0.714f
C3103 m1_4468_94364# m2_4468_94364# 12.9f
C3104 xaa0.xa5.MN2.G xaa6.xc.XA7.MN0.D 0.12f
C3105 xaa6.xc.XA1.MN0.G xaa6.xc.XA7.MN1.G 0.412f
C3106 a_32284_58030# xaa6.xe.XA7.MP1.G 3.8e-19
C3107 a_27244_57678# a_28612_57678# 8.89e-19
C3108 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MP1.G 0.313f
C3109 xaa6.xe.XA1.MN0.G a_34804_57678# 0.00417f
C3110 xaa6.xf.XA7.MN1.D a_33652_57678# 0.0877f
C3111 AVDD a_n908_55566# 0.00171f
C3112 xaa6.xe.XA1.MN0.G a_31132_54158# 0.00118f
C3113 xaa6.xe.XA7.MN1.D a_32284_54158# 0.0747f
C3114 xaa6.xe.XA6.MN0.G xaa6.xf.XA6.MN0.G 0.00435f
C3115 a_2948_74698# li_4468_75004# 8.34e-20
C3116 xaa1.xa4.M0.D li_4468_74044# 23f
C3117 AVDD a_34804_52750# 0.00535f
C3118 xaa1.xa4.M0.D m3_4788_98364# 0.0138f
C3119 xaa4.xa1.M6.D xaa4.xa1.M5.D 0.0488f
C3120 li_4468_106684# li_4468_105884# 39.3f
C3121 a_28612_64622# xaa5.xb1.MN1.G 2.54e-19
C3122 xaa3.xa3a.MN0.D a_5844_58494# 0.0536f
C3123 AVDD a_31132_57678# 0.00163f
C3124 xaa6.xg.XA7.MP1.G a_37324_55918# 0.0292f
C3125 xaa0.xa5.MP1.D a_244_55918# 0.0494f
C3126 AVDD a_27244_54158# 0.387f
C3127 a_4692_55150# a_4308_53678# 0.00374f
C3128 a_10092_55038# a_10092_54510# 0.00702f
C3129 xaa6.xg.XA5.MN0.G a_37324_54158# 1.28e-19
C3130 xaa1.xa4.M0.D m3_37668_114844# 0.074f
C3131 a_37324_56270# m1_37504_55818# 0.00413f
C3132 li_4468_93404# m1_4468_93404# 23f
C3133 xaa5.xb1.MN1.D a_29764_61454# 0.127f
C3134 AVDD a_28612_61454# 0.352f
C3135 a_n940_74698# a_n508_74698# 0.00813f
C3136 m2_4468_115484# m3_37748_115804# 0.0138f
C3137 xaa6.xg.XA7.MN1.G xaa6.xg.XA7.MN2.D 0.0148f
C3138 xaa6.xg.XA7.MP1.G xaa6.xg.XA7.MN0.G 0.0605f
C3139 xaa6.xe.XA7.MP1.G a_31132_56974# 2.35e-19
C3140 xaa6.xe.XA7.MN1.G a_32284_56974# 0.0035f
C3141 a_n908_56974# a_244_56974# 0.00133f
C3142 xaa6.xc.XA7.MN1.G a_27244_56622# 0.0769f
C3143 xaa6.xc.XA7.MP1.G a_26092_56622# 0.0692f
C3144 AVDD a_244_54862# 0.386f
C3145 a_36172_55566# a_37324_55566# 0.00133f
C3146 xaa6.xf.XA1.MN0.G a_34804_52750# 0.00159f
C3147 xaa6.xd.XA7.MN1.G a_29764_53102# 7.28e-19
C3148 xaa6.xc.XA6.MN0.G a_27244_54862# 0.0725f
C3149 a_29764_53806# a_29764_53454# 0.0109f
C3150 xaa1.xa4.M0.D m3_37748_81244# 0.111f
C3151 li_4468_89564# li_4468_89404# 7.91f
C3152 xaa0.xa6.MN0.D xaa1.xa1.M8.D 4.21e-19
C3153 xaa5.xb1.MN1.G xaa5.xb2_0.MN0.D 0.0438f
C3154 xaa5.xa3.xb2_0.G a_27244_62158# 0.00147f
C3155 AVDD xaa0.xa6.MN0.D 1.43f
C3156 m1_4468_70364# m1_4468_70204# 11.3f
C3157 IBPSR_1U xaa4.xa1.M8.D 0.0166f
C3158 PWRUP_1V8 a_n908_55918# 3.01e-19
C3159 a_32284_58030# xaa6.xe.XA7.MN1.G 3.89e-19
C3160 xaa0.xa5.MN2.G xaa6.xc.XA7.MP1.G 0.193f
C3161 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MN1.G 0.467f
C3162 xaa6.xe.XA1.MN0.G a_33652_57678# 0.0258f
C3163 AVDD xaa0.xa1.MN0.G 1.23f
C3164 xaa6.xe.XA7.MN1.D a_31132_54158# 0.066f
C3165 xaa6.xg.XA6.MP0.D a_37324_55918# 0.00176f
C3166 a_31132_56270# a_31132_55918# 0.0109f
C3167 xaa6.xd.XA1.MN0.G a_32284_54158# 1.11e-19
C3168 a_2948_74698# li_4468_75164# 3.68e-19
C3169 xaa4.xa4.M0.D xaa4.xa1.M2.D 4.85e-19
C3170 xaa6.xc.XA7.MN1.G a_28612_54510# 7.1e-20
C3171 xaa6.xc.XA7.MP1.G a_27244_54510# 0.0969f
C3172 AVDD a_33652_52750# 0.447f
C3173 xaa1.xa4.M0.D m3_4628_98364# 0.0276f
C3174 a_32284_54510# a_32284_54158# 0.0109f
C3175 xaa1.xa4.M0.G xaa3.xa8.MP0.D 0.062f
C3176 xaa1.xa3.D xaa4.xa2.M0.G 0.746f
C3177 a_4692_63774# a_5844_63774# 0.00133f
C3178 a_4692_64126# xaa3.xa7.MN0.D 4.14e-19
C3179 li_4468_71324# m1_4468_71324# 23f
C3180 xaa3.xa3a.MN0.D a_4692_58494# 0.0583f
C3181 a_28612_60750# a_29764_60750# 0.00133f
C3182 AVDD a_29764_57678# 0.00163f
C3183 m2_4468_102044# m3_37748_102364# 0.0138f
C3184 xaa1.xa4.M0.D li_4468_108604# 23f
C3185 xaa6.xd.XA7.MN1.G xaa6.xd.XA5.MN0.G 0.0911f
C3186 xaa0.xa5.MN2.G a_n908_53806# 4.05e-20
C3187 xaa6.xg.XA7.MN1.G a_37324_55918# 0.00718f
C3188 xaa6.xg.XA7.MP1.G a_36172_55918# 0.0294f
C3189 AVDD a_26092_54158# 0.00164f
C3190 xaa4.xa2.M0.D xaa4.xa1.M3.D 0.00219f
C3191 a_37324_55214# xaa6.xg.XA4.MN0.G 0.0658f
C3192 a_31132_55214# a_31132_54862# 0.0109f
C3193 xaa6.xg.XA5.MN0.G a_36172_54158# 1.95e-19
C3194 xaa1.xa4.M0.D m3_4788_115644# 0.0138f
C3195 xbb1.xa3.M3.D xbb1.xa3.M2.D 0.0488f
C3196 a_29764_52750# a_31132_52750# 8.89e-19
C3197 a_37324_56270# m1_37504_57930# 1.49e-19
C3198 li_4468_73084# li_4468_72284# 39.3f
C3199 xaa5.xb1.MN1.D a_28612_61454# 0.0685f
C3200 a_n908_61510# xaa1.xa1.M6.D 5.84e-19
C3201 xaa3.xa1b.MN0.D xaa0.xa5.MN2.G 5.43e-19
C3202 AVDD a_27244_61454# 0.382f
C3203 m2_4468_115484# m3_37668_115804# 0.0138f
C3204 xaa6.xg.XA7.MN1.G xaa6.xg.XA7.MN0.G 0.041f
C3205 xaa6.xe.XA7.MN1.G a_31132_56974# 0.00922f
C3206 xaa6.xc.XA7.MN1.G a_26092_56622# 0.0111f
C3207 PWRUP_1V8 a_36172_55566# 0.00493f
C3208 AVDD a_n908_54862# 0.00171f
C3209 xaa1.xa4.M0.D m1_4468_72284# 56.4f
C3210 a_2948_74698# m1_4468_74204# 5.04e-19
C3211 xaa6.xc.XA5.MN0.G xaa6.xc.XA4.MP0.D 0.0618f
C3212 xaa0.xa5.MN2.G a_4308_51566# 9.74e-19
C3213 xaa6.xf.XA7.MN1.D a_34804_52750# 6.12e-22
C3214 xaa6.xd.XA7.MN1.G a_28612_53102# 0.00893f
C3215 xaa6.xd.XA7.MP1.G a_29764_53102# 1.1e-19
C3216 xaa6.xc.XA6.MN0.G a_26092_54862# 0.0658f
C3217 a_36172_53806# xaa6.xg.XA1.MN0.D 0.00176f
C3218 xaa1.xa4.M0.D m3_37668_81244# 0.074f
C3219 li_4468_116444# m1_4468_116444# 23f
C3220 a_27244_63214# a_28612_63214# 8.89e-19
C3221 xaa5.xa3.xb2_0.G a_26092_62158# 0.0767f
C3222 IBPSR_1U xaa1.xa2.M0.D 0.026f
C3223 xaa4.xa2.M0.G a_29764_62158# 3.48e-19
C3224 AVDD a_n908_63622# 7.8e-20
C3225 m1_4468_95324# m2_4468_95324# 12.9f
C3226 a_31132_58030# xaa6.xe.XA7.MN1.G 8.24e-19
C3227 a_26092_57678# a_27244_57678# 0.00133f
C3228 xaa0.xa5.MN2.G xaa6.xc.XA7.MN1.G 0.0632f
C3229 xaa6.xe.XA1.MN0.G a_32284_57678# 0.00249f
C3230 AVDD a_244_55918# 0.364f
C3231 m2_4468_88604# m3_37748_88924# 0.0138f
C3232 xaa6.xd.XA1.MN0.G a_31132_54158# 0.00207f
C3233 xaa6.xe.XA7.MP1.G xaa6.xe.XA3.MP0.D 0.0712f
C3234 a_2948_74698# li_4468_75964# 1.04e-19
C3235 xaa1.xa4.M0.D li_4468_75004# 23f
C3236 PWRUP_1V8 a_29764_52750# 4.95e-20
C3237 xaa6.xc.XA7.MN1.G a_27244_54510# 0.0057f
C3238 xaa6.xc.XA7.MP1.G a_26092_54510# 0.0278f
C3239 xaa6.xd.XA6.MN0.G xaa6.xe.XA6.MN0.G 0.00435f
C3240 a_37324_56270# xaa6.xg.XA6.MN0.G 0.0658f
C3241 AVDD a_32284_52750# 0.449f
C3242 xaa1.xa4.M0.D m3_37748_98524# 0.111f
C3243 li_4468_106844# li_4468_106684# 7.91f
C3244 xaa1.xa4.M0.G xaa3.xa7.MN0.D 0.347f
C3245 xaa3.xa9.MN0.D a_5844_63774# 0.00224f
C3246 xaa1.xb1.M0.D a_640_59750# 0.00155f
C3247 xaa0.xa2a.MN0.D xaa0.xa5.MN2.G 0.00172f
C3248 PWRUP_1V8 a_26092_57678# 0.00459f
C3249 AVDD a_28612_57678# 0.384f
C3250 m2_4468_102044# m3_37668_102364# 0.0138f
C3251 xaa6.xd.XA7.MN1.G xaa6.xc.XA5.MN0.G 1.74e-19
C3252 xaa6.xd.XA7.MP1.G xaa6.xd.XA5.MN0.G 0.397f
C3253 xaa6.xg.XA7.MN1.D a_37324_55566# 0.00147f
C3254 xaa6.xg.XA7.MN1.G a_36172_55918# 7.37e-19
C3255 AVDD xaa4.xa1.M5.D 0.00415f
C3256 xaa4.xa2.M0.D xaa4.xa1.M4.D 0.00265f
C3257 xaa6.xg.XA4.MP0.D a_37324_54862# 0.00176f
C3258 a_36172_55214# xaa6.xg.XA4.MN0.G 0.0674f
C3259 xaa1.xa4.M0.D m3_4628_115644# 0.0276f
C3260 xaa1.xa1.M7.D PWRUP_1V8 0.0119f
C3261 IBPSR_1U xaa0.xa5.MN2.G 0.0278f
C3262 AVDD a_26092_61454# 0.00164f
C3263 a_n940_74698# xbb0.xa1.XA1.N 0.104f
C3264 a_26092_57326# xaa6.xc.XA7.MN2.D 0.00176f
C3265 PWRUP_1V8 a_34804_55566# 0.00493f
C3266 AVDD a_37324_55566# 0.383f
C3267 m2_4468_75164# m3_37748_75484# 0.0138f
C3268 xaa1.xa4.M0.D m1_4468_73244# 67.7f
C3269 a_2948_74698# m1_4468_75164# 0.00161f
C3270 a_34804_55566# a_36172_55566# 8.89e-19
C3271 xaa6.xf.XA7.MN1.G a_34804_53454# 0.015f
C3272 xaa6.xc.XA5.MN0.G xaa6.xc.XA4.MN0.D 0.126f
C3273 xaa6.xf.XA7.MN1.D a_33652_52750# 3.67e-21
C3274 xaa6.xf.XA6.MN0.G a_34804_55214# 0.0658f
C3275 a_28612_53806# a_28612_53454# 0.0109f
C3276 xaa1.xa4.M0.D m3_4788_82044# 0.0138f
C3277 li_4468_90364# li_4468_89564# 39.3f
C3278 a_n908_63270# xaa1.xa2.M0.D 5.02e-20
C3279 xaa4.xa2.M0.G a_28612_62158# 0.0362f
C3280 AVDD a_5844_63774# 0.384f
C3281 m1_4468_71164# m1_4468_70364# 56.4f
C3282 xaa6.xd.XA1.MN0.G a_33652_57678# 2.93e-19
C3283 PWRUP_1V8 a_37324_56622# 0.0674f
C3284 xaa6.xe.XA7.MN1.D a_32284_57678# 0.0893f
C3285 xaa6.xe.XA1.MN0.G a_31132_57678# 1.35e-19
C3286 AVDD a_n908_55918# 0.00164f
C3287 m2_4468_88604# m3_37668_88924# 0.0138f
C3288 a_29764_56270# a_29764_55918# 0.0109f
C3289 xaa6.xg.XA6.MN0.D a_36172_55918# 0.00176f
C3290 xaa6.xg.XA7.MP1.G a_37324_54862# 0.097f
C3291 xaa6.xd.XA1.MN0.G a_29764_54158# 0.00268f
C3292 xaa6.xe.XA7.MP1.G xaa6.xe.XA3.MN0.D 0.0472f
C3293 xaa6.xe.XA7.MN1.G xaa6.xe.XA3.MP0.D 0.00252f
C3294 a_2948_74698# li_4468_76124# 3.68e-19
C3295 xaa6.xc.XA7.MN1.G a_26092_54510# 0.082f
C3296 a_36172_56270# xaa6.xg.XA6.MN0.G 0.0674f
C3297 AVDD a_31132_52750# 0.00535f
C3298 xaa1.xa4.M0.D m3_37668_98524# 0.074f
C3299 xaa4.xa1.M7.D xaa4.xa1.M6.D 0.0488f
C3300 a_31132_54510# a_31132_54158# 0.0109f
C3301 xaa6.xg.XA3.MP0.D a_37324_54158# 0.00176f
C3302 xaa1.xa4.M0.G xaa0.xa6.MN0.D 0.25f
C3303 a_5844_64126# a_5844_63774# 0.0109f
C3304 xaa3.xa9.MN0.D a_4692_63774# 0.00224f
C3305 li_4468_72124# m1_4468_72124# 23f
C3306 a_27244_60750# a_28612_60750# 8.89e-19
C3307 PWRUP_1V8 xaa6.xg.XA7.MN1.D 0.16f
C3308 AVDD a_27244_57678# 0.384f
C3309 xaa6.xg.XA7.MN1.D a_36172_55566# 0.00699f
C3310 xaa1.xa4.M0.D li_4468_109564# 23f
C3311 xaa0.xa5.MN2.G xaa0.xa1.MN0.D 9.89e-20
C3312 xaa6.xf.XA1.MN0.G a_37324_55566# 1.11e-19
C3313 AVDD xaa4.xa1.M6.D 0.00415f
C3314 a_36172_55214# a_37324_55214# 0.00133f
C3315 a_29764_55214# a_29764_54862# 0.0109f
C3316 xaa1.xa4.M0.D m3_37748_115804# 0.111f
C3317 xaa3.xa4.MN0.D li_4980_61284# 7.61e-20
C3318 a_37324_53102# a_37324_52750# 0.0109f
C3319 a_28612_52750# a_29764_52750# 0.00133f
C3320 xaa1.xa3.D m3_4788_69564# 0.0138f
C3321 li_4468_73244# li_4468_73084# 7.91f
C3322 li_4468_94364# m1_4468_94364# 23f
C3323 a_29764_61806# a_29764_61454# 0.0109f
C3324 xaa1.xa1.M8.D PWRUP_1V8 0.25f
C3325 AVDD PWRUP_1V8 15.3f
C3326 xaa6.xf.XA7.MN0.D xaa6.xf.XA7.MN2.D 0.0618f
C3327 xaa0.xa5.MN2.G xaa0.xa1.MN2.S 8.83e-19
C3328 xaa6.xd.XA7.MN0.D a_29764_56974# 0.00297f
C3329 AVDD a_36172_55566# 0.00151f
C3330 m2_4468_75164# m3_37668_75484# 0.0138f
C3331 xaa6.xf.XA7.MP1.G a_34804_53454# 2.78e-19
C3332 xaa6.xf.XA7.MN1.G a_33652_53454# 0.101f
C3333 xaa1.xa4.M0.D m1_4468_74204# 67.7f
C3334 a_2948_74698# m1_4468_76124# 0.00161f
C3335 xaa6.xf.XA6.MN0.G a_33652_55214# 0.0827f
C3336 a_34804_53806# xaa6.xf.XA1.MN0.D 0.00176f
C3337 xaa1.xa4.M0.D m3_4628_82044# 0.0276f
C3338 xaa0.xa6.MN0.D a_n908_61510# 8.05e-19
C3339 xaa5.xa3.xb2_0.G xaa5.xb2_1.MN0.D 0.0025f
C3340 a_26092_63214# a_27244_63214# 0.00133f
C3341 xaa5.xb1.MN1.G a_29764_62158# 0.00585f
C3342 xaa4.xa2.M0.G a_27244_62158# 6.34e-19
C3343 AVDD a_4692_63774# 0.00171f
C3344 m1_4468_96284# m2_4468_96284# 12.9f
C3345 xaa6.xd.XA1.MN0.G a_32284_57678# 0.021f
C3346 PWRUP_1V8 a_36172_56622# 0.0777f
C3347 xaa4.xa2.M0.G a_10092_55566# 0.00391f
C3348 xaa6.xe.XA7.MN1.D a_31132_57678# 0.132f
C3349 AVDD xaa0.xa5.MP1.D 0.191f
C3350 xaa6.xg.XA7.MP1.G a_36172_54862# 0.029f
C3351 xaa6.xg.XA7.MN1.G a_37324_54862# 0.00639f
C3352 xaa6.xd.XA7.MN1.D a_29764_54158# 0.0676f
C3353 xaa6.xd.XA1.MN0.G a_28612_54158# 1.35e-19
C3354 xaa6.xe.XA7.MN1.G xaa6.xe.XA3.MN0.D 0.0288f
C3355 a_2948_74698# li_4468_76924# 1.04e-19
C3356 xaa1.xa4.M0.D li_4468_75964# 23f
C3357 xaa6.xc.XA6.MN0.G xaa6.xd.XA6.MN0.G 0.00435f
C3358 AVDD a_29764_52750# 0.00535f
C3359 xaa1.xa4.M0.D m3_4788_99324# 0.0138f
C3360 a_10092_54510# xaa4.xa1.M3.D 1.21e-19
C3361 li_4468_107644# li_4468_106844# 39.3f
C3362 xaa1.xa4.M0.G a_n908_63622# 0.0733f
C3363 PWRUP_1V8 xaa6.xf.XA1.MN0.G 0.456f
C3364 AVDD a_26092_57678# 0.00171f
C3365 xaa6.xf.XA1.MN0.G a_36172_55566# 0.00205f
C3366 a_33652_57326# xaa6.xf.XA6.MN0.G 5e-20
C3367 AVDD a_11712_54334# 0.424f
C3368 xaa6.xf.XA5.MN0.G a_34804_54158# 1.95e-19
C3369 xaa6.xg.XA4.MN0.D a_36172_54862# 0.00176f
C3370 xaa1.xa4.M0.D m3_37668_115804# 0.074f
C3371 xaa3.xa4.MN0.D li_4836_61284# 4.62e-19
C3372 xaa1.xa3.D m3_4628_69564# 0.0276f
C3373 xaa5.xb1.MN1.D PWRUP_1V8 0.0542f
C3374 xaa1.xa1.M8.D xaa1.xa1.M7.D 0.063f
C3375 a_36172_57326# a_37324_57326# 0.00133f
C3376 xaa6.xg.XA7.MN1.D a_37324_56622# 0.0232f
C3377 xaa6.xf.XA7.MN1.G xaa6.xf.XA7.MN2.D 0.0148f
C3378 xaa6.xd.XA7.MN1.G a_29764_56974# 0.00922f
C3379 xaa6.xd.XA7.MN0.D a_28612_56974# 0.016f
C3380 AVDD a_34804_55566# 0.00151f
C3381 xaa6.xf.XA7.MP1.G a_33652_53454# 1.07e-19
C3382 xaa6.xf.XA7.MN1.G a_32284_53454# 7.1e-20
C3383 xaa1.xa4.M0.D m1_4468_75164# 67.7f
C3384 a_2948_74698# m1_4468_77084# 5.67e-19
C3385 a_33652_55566# a_34804_55566# 0.00133f
C3386 xaa6.xe.XA1.MN0.G a_32284_52750# 0.00177f
C3387 a_27244_53806# a_27244_53454# 0.0109f
C3388 xaa1.xa4.M0.D m3_37748_82204# 0.111f
C3389 li_4468_117404# m1_4468_117404# 23f
C3390 li_4468_90524# li_4468_90364# 7.91f
C3391 xaa1.xa3.D xaa0.xa2a.MN0.D 0.0185f
C3392 xaa5.xa3.xb2_0.G xaa5.xa3.xb1_0.D 0.294f
C3393 IBPSR_1U xaa1.xa2.M1.D 0.026f
C3394 xaa5.xb1.MN1.G a_28612_62158# 9.6e-19
C3395 AVDD xaa3.xa9.MN0.D 0.176f
C3396 m1_4468_71324# m1_4468_71164# 11.3f
C3397 a_29764_58030# xaa6.xd.XA7.MN1.G 0.00227f
C3398 xaa6.xd.XA1.MN0.G a_31132_57678# 0.00739f
C3399 PWRUP_1V8 a_34804_56622# 0.0796f
C3400 a_37324_58030# a_37324_57678# 0.0109f
C3401 AVDD a_37324_56622# 0.364f
C3402 a_28612_56270# a_28612_55918# 0.0109f
C3403 xaa6.xf.XA6.MN0.D a_34804_55918# 0.00176f
C3404 xaa6.xg.XA7.MN1.G a_36172_54862# 1.25e-19
C3405 xaa6.xd.XA7.MN1.D a_28612_54158# 0.0731f
C3406 xaa6.xc.XA1.MN0.G a_29764_54158# 1.11e-19
C3407 a_2948_74698# li_4468_77084# 1.28e-19
C3408 PWRUP_1V8 a_26092_52750# 4.2e-19
C3409 a_34804_56270# xaa6.xf.XA6.MN0.G 0.0661f
C3410 AVDD a_28612_52750# 0.447f
C3411 xaa1.xa4.M0.D m3_4628_99324# 0.0276f
C3412 a_10092_54510# xaa4.xa1.M4.D 1.81e-19
C3413 a_29764_54510# a_29764_54158# 0.0109f
C3414 xaa6.xg.XA3.MN0.D a_36172_54158# 0.00176f
C3415 xaa6.xg.XA3.MN1.G a_37324_54158# 0.0676f
C3416 xaa1.xa3.D IBPSR_1U 0.00876f
C3417 a_4692_64126# a_4692_63774# 0.0109f
C3418 xaa1.xa4.M0.G a_5844_63774# 0.0921f
C3419 a_n908_64150# a_n908_63622# 0.00702f
C3420 a_5844_64126# xaa3.xa9.MN0.D 0.0215f
C3421 li_4468_72284# m1_4468_72284# 23f
C3422 a_640_60278# a_640_59750# 0.00702f
C3423 PWRUP_1V8 xaa6.xf.XA7.MN1.D 0.161f
C3424 xaa1.xa1.M0.D a_n908_59750# 0.00155f
C3425 a_26092_60750# a_27244_60750# 0.00133f
C3426 CK xaa6.xg.XA7.MN0.D 6.8e-19
C3427 AVDD xaa6.xg.XA7.MN1.D 1.86f
C3428 xaa6.xf.XA7.MN1.G a_34804_55918# 7.37e-19
C3429 PWRUP_1V8 a_36172_54510# 0.00467f
C3430 xaa1.xa4.M0.D li_4468_110524# 23f
C3431 xaa0.xa5.MN2.G a_n908_54158# 4.05e-20
C3432 xaa6.xf.XA1.MN0.G a_34804_55566# 0.00217f
C3433 xaa6.xc.XA7.MN1.G xaa6.xd.XA5.MN0.G 1.74e-19
C3434 xaa6.xc.XA7.MP1.G xaa6.xc.XA5.MN0.G 0.397f
C3435 a_36172_56622# a_37324_56622# 0.00133f
C3436 AVDD xaa4.xa1.M7.D 0.00415f
C3437 xaa6.xf.XA5.MN0.G a_33652_54158# 1.28e-19
C3438 a_34804_55214# a_36172_55214# 8.89e-19
C3439 a_28612_55214# a_28612_54862# 0.0109f
C3440 xaa1.xa4.M0.D m3_4788_116604# 0.0138f
C3441 a_36172_53102# a_36172_52750# 0.0109f
C3442 a_27244_52750# a_28612_52750# 8.89e-19
C3443 xaa1.xa3.D m3_37748_69724# 0.111f
C3444 li_4468_74044# li_4468_73244# 39.3f
C3445 a_640_61510# PWRUP_1V8 0.069f
C3446 a_28612_61806# a_28612_61454# 0.0109f
C3447 AVDD xaa1.xa1.M8.D 2.27f
C3448 m2_4468_116444# m3_37748_116764# 0.0138f
C3449 xaa6.xg.XA7.MN1.D a_36172_56622# 0.0377f
C3450 xaa0.xa5.MN2.G a_n908_55214# 2.3e-19
C3451 PWRUP_1V8 a_31132_55566# 0.00493f
C3452 xaa6.xd.XA7.MP1.G a_29764_56974# 2.35e-19
C3453 xaa6.xd.XA7.MN1.G a_28612_56974# 0.0035f
C3454 AVDD a_33652_55566# 0.383f
C3455 xaa1.xa4.M0.D m1_4468_76124# 67.7f
C3456 xaa6.xe.XA7.MN1.D a_32284_52750# 3.67e-21
C3457 xaa6.xe.XA1.MN0.G a_31132_52750# 0.00263f
C3458 xaa6.xe.XA6.MN0.G a_32284_55214# 0.0811f
C3459 xaa4.xa1.M5.D a_10092_52750# 8.62e-20
C3460 xaa1.xa4.M0.D m3_37668_82204# 0.074f
C3461 xaa5.xa3.xb2_0.G xaa5.xa4.MN0.D 0.011f
C3462 a_n908_63270# xaa1.xa2.M1.D 6.46e-20
C3463 xaa5.xa3.xb1_0.G a_26092_62158# 0.00208f
C3464 AVDD a_5844_64126# 0.351f
C3465 m1_4468_97244# m2_4468_97244# 12.9f
C3466 a_28612_58030# xaa6.xd.XA7.MN1.G 1.55e-20
C3467 xaa6.xd.XA1.MN0.G a_29764_57678# 0.00219f
C3468 PWRUP_1V8 a_33652_56622# 0.0658f
C3469 xaa6.xf.XA1.MN0.G xaa6.xg.XA7.MN1.D 0.147f
C3470 AVDD a_36172_56622# 0.00151f
C3471 xaa6.xc.XA1.MN0.G a_28612_54158# 0.00209f
C3472 a_2948_74698# li_4468_77884# 1.76e-20
C3473 xaa1.xa4.M0.D li_4468_76924# 23f
C3474 PWRUP_1V8 a_11712_52750# 0.00173f
C3475 xaa6.xg.XA7.MN1.D a_37324_54510# 0.0836f
C3476 a_33652_56270# xaa6.xf.XA6.MN0.G 0.0735f
C3477 AVDD a_27244_52750# 0.449f
C3478 xaa1.xa4.M0.D m3_37748_99484# 0.111f
C3479 xaa6.xg.XA3.MN1.G a_36172_54158# 0.08f
C3480 li_4468_107804# li_4468_107644# 7.91f
C3481 xaa1.xa3.D a_n908_63270# 0.00678f
C3482 a_4692_64126# xaa3.xa9.MN0.D 0.0215f
C3483 xaa1.xa4.M0.G a_4692_63774# 0.0951f
C3484 PWRUP_1V8 xaa6.xe.XA1.MN0.G 0.209f
C3485 CK xaa6.xg.XA7.MP1.G 0.00168f
C3486 AVDD xaa6.xf.XA1.MN0.G 0.757f
C3487 m2_4468_103004# m3_37748_103324# 0.0138f
C3488 xaa6.xf.XA7.MN1.G a_33652_55918# 0.00733f
C3489 xaa6.xf.XA7.MP1.G a_34804_55918# 0.0294f
C3490 PWRUP_1V8 a_34804_54510# 0.00467f
C3491 xaa6.xf.XA7.MN1.D a_34804_55566# 0.00699f
C3492 xaa6.xc.XA7.MN1.G xaa6.xc.XA5.MN0.G 0.0911f
C3493 a_32284_57326# xaa6.xe.XA6.MN0.G 5e-20
C3494 xaa6.xf.XA1.MN0.G a_33652_55566# 1.35e-19
C3495 AVDD a_37324_54510# 0.362f
C3496 xaa1.xa4.M0.D m3_4628_116604# 0.0276f
C3497 xaa1.xa3.D m3_37668_69724# 0.074f
C3498 li_4468_95324# m1_4468_95324# 23f
C3499 a_n908_61510# PWRUP_1V8 0.00637f
C3500 AVDD xaa5.xb1.MN1.D 0.636f
C3501 m2_4468_116444# m3_37668_116764# 0.0138f
C3502 a_34804_57326# a_36172_57326# 8.89e-19
C3503 PWRUP_1V8 a_29764_55566# 0.00493f
C3504 xaa6.xf.XA1.MN0.G a_36172_56622# 0.00133f
C3505 xaa6.xd.XA7.MP1.G a_28612_56974# 0.0291f
C3506 AVDD a_32284_55566# 0.383f
C3507 xaa6.xc.XA7.MP1.G a_26092_53102# 1.1e-19
C3508 xaa6.xc.XA7.MN1.G a_27244_53102# 0.00893f
C3509 xaa1.xa4.M0.D m1_4468_77084# 67.7f
C3510 a_32284_55566# a_33652_55566# 8.89e-19
C3511 xaa6.xe.XA7.MN1.D a_31132_52750# 6.12e-22
C3512 xaa6.xe.XA6.MN0.G a_31132_55214# 0.0674f
C3513 xaa4.xa1.M6.D a_10092_52750# 6.46e-20
C3514 a_26092_53806# a_26092_53454# 0.0109f
C3515 a_11712_54334# a_11712_52750# 0.00223f
C3516 xaa1.xa4.M0.D m3_4788_83004# 0.0138f
C3517 li_4468_91324# li_4468_90524# 39.3f
C3518 xaa4.xa2.M0.G xaa5.xb2_1.MN0.D 0.174f
C3519 xaa5.xa3.xb2_0.G a_29764_62510# 1.93e-19
C3520 AVDD a_4692_64126# 0.00623f
C3521 m1_4468_72124# m1_4468_71324# 56.4f
C3522 xaa6.xd.XA1.MN0.G a_28612_57678# 1.35e-19
C3523 a_28612_58030# xaa6.xd.XA7.MP1.G 3.8e-19
C3524 xaa6.xd.XA7.MN1.D a_29764_57678# 0.134f
C3525 PWRUP_1V8 a_32284_56622# 0.0674f
C3526 a_36172_58030# a_36172_57678# 0.0109f
C3527 xaa6.xf.XA7.MN1.D xaa6.xg.XA7.MN1.D 0.00642f
C3528 AVDD a_34804_56622# 0.00151f
C3529 m2_4468_89564# m3_37748_89884# 0.0138f
C3530 a_27244_56270# a_27244_55918# 0.0109f
C3531 xaa6.xf.XA6.MP0.D a_33652_55918# 0.00176f
C3532 xaa6.xd.XA7.MN1.G xaa6.xd.XA3.MN0.D 0.0288f
C3533 xaa6.xf.XA1.MN0.G a_37324_54510# 1.11e-19
C3534 xaa6.xc.XA1.MN0.G a_27244_54158# 0.00329f
C3535 PWRUP_1V8 a_10092_52750# 0.00152f
C3536 xaa6.xg.XA7.MN1.D a_36172_54510# 0.0736f
C3537 AVDD a_26092_52750# 0.00543f
C3538 xaa1.xa4.M0.D m3_37668_99484# 0.074f
C3539 a_28612_54510# a_28612_54158# 0.0109f
C3540 a_4692_64126# a_5844_64126# 0.00133f
C3541 xaa1.xa4.M0.G xaa3.xa9.MN0.D 0.17f
C3542 PWRUP_1V8 xaa6.xe.XA7.MN1.D 0.16f
C3543 CK xaa6.xg.XA7.MN1.G 0.293f
C3544 xaa1.xa1.M1.D a_n908_59750# 5.84e-19
C3545 AVDD xaa6.xf.XA7.MN1.D 1.86f
C3546 m2_4468_103004# m3_37668_103324# 0.0138f
C3547 xaa6.xf.XA7.MN1.G a_32284_55918# 7.1e-20
C3548 xaa6.xf.XA7.MP1.G a_33652_55918# 0.0292f
C3549 xaa1.xa4.M0.D li_4468_111484# 23f
C3550 xaa0.xa5.MN2.G a_n908_54510# 1.97e-19
C3551 xaa6.xf.XA7.MN1.D a_33652_55566# 0.00147f
C3552 xaa6.xe.XA1.MN0.G a_34804_55566# 1.02e-19
C3553 a_34804_56622# a_36172_56622# 8.89e-19
C3554 AVDD a_36172_54510# 0.00151f
C3555 xaa6.xf.XA4.MN0.D a_34804_54862# 0.00176f
C3556 a_33652_55214# a_34804_55214# 0.00133f
C3557 a_27244_55214# a_27244_54862# 0.0109f
C3558 xaa1.xa4.M0.D m3_37748_116764# 0.111f
C3559 a_4692_60782# li_4980_61284# 2e-19
C3560 xaa6.xe.XA5.MN0.G a_32284_54158# 1.28e-19
C3561 a_34804_53102# a_34804_52750# 0.0109f
C3562 a_26092_52750# a_27244_52750# 0.00133f
C3563 xaa1.xa3.D m3_4788_70524# 0.0138f
C3564 li_4468_74204# li_4468_74044# 7.91f
C3565 a_29764_61806# PWRUP_1V8 4.95e-20
C3566 a_640_61510# xaa1.xa1.M8.D 0.0124f
C3567 a_n908_61510# xaa1.xa1.M7.D 0.00155f
C3568 a_27244_61806# a_27244_61454# 0.0109f
C3569 AVDD a_640_61510# 0.333f
C3570 xaa6.xe.XA7.MN0.D xaa6.xe.XA7.MN2.D 0.0618f
C3571 xaa6.xf.XA1.MN0.G a_34804_56622# 0.00134f
C3572 AVDD a_31132_55566# 0.00151f
C3573 m2_4468_76124# m3_37748_76444# 0.0138f
C3574 xaa6.xc.XA7.MN1.G a_26092_53102# 7.44e-19
C3575 xaa3.xa1b.MN0.D li_4980_56708# 3.78e-19
C3576 xaa1.xa4.M0.D m1_4468_78044# 67.7f
C3577 xaa6.xe.XA7.MN1.G a_33652_53454# 7.1e-20
C3578 xaa6.xe.XA7.MP1.G a_32284_53454# 1.07e-19
C3579 a_31132_53806# xaa6.xe.XA1.MN0.D 0.00176f
C3580 xaa1.xa4.M0.D m3_4628_83004# 0.0276f
C3581 xaa4.xa2.M0.G xaa5.xa3.xb1_0.D 0.012f
C3582 xaa5.xa3.xb2_0.G a_28612_62510# 8.96e-19
C3583 a_4692_62366# a_5844_62366# 0.00133f
C3584 AVDD xaa1.xa4.M0.G 2.45f
C3585 m1_4468_98204# m2_4468_98204# 12.9f
C3586 xaa6.xd.XA7.MN1.D a_28612_57678# 0.0877f
C3587 xaa6.xf.XA7.MN1.D xaa6.xf.XA1.MN0.G 0.0167f
C3588 xaa6.xc.XA1.MN0.G a_29764_57678# 0.00417f
C3589 PWRUP_1V8 a_31132_56622# 0.0777f
C3590 xaa3.xa1b.MN0.D a_5844_55150# 1.28e-19
C3591 xaa6.xe.XA1.MN0.G xaa6.xg.XA7.MN1.D 2.06e-19
C3592 AVDD a_33652_56622# 0.365f
C3593 m2_4468_89564# m3_37668_89884# 0.0138f
C3594 xaa6.xd.XA7.MN1.G xaa6.xd.XA3.MP0.D 0.00252f
C3595 xaa6.xd.XA7.MP1.G xaa6.xd.XA3.MN0.D 0.0472f
C3596 xaa6.xf.XA1.MN0.G a_36172_54510# 0.00193f
C3597 xaa6.xc.XA7.MN1.D a_27244_54158# 0.0747f
C3598 xaa6.xc.XA1.MN0.G a_26092_54158# 0.00118f
C3599 a_5844_55854# a_5844_55502# 0.0109f
C3600 xaa1.xa4.M0.D li_4468_77884# 23f
C3601 xaa6.xf.XA7.MN1.G a_34804_54862# 0.0708f
C3602 a_36172_56270# a_37324_56270# 0.00133f
C3603 a_32284_56270# xaa6.xe.XA6.MN0.G 0.0719f
C3604 AVDD a_11712_52750# 0.395f
C3605 xaa1.xa4.M0.D m3_4788_100284# 0.0138f
C3606 a_36172_54510# a_37324_54510# 0.00133f
C3607 xaa6.xf.XA3.MN0.D a_34804_54158# 0.00176f
C3608 li_4468_108604# li_4468_107804# 39.3f
C3609 xaa1.xa4.M0.G a_5844_64126# 0.069f
C3610 li_4468_73244# m1_4468_73244# 23f
C3611 PWRUP_1V8 xaa6.xd.XA1.MN0.G 0.537f
C3612 AVDD xaa6.xe.XA1.MN0.G 3.52f
C3613 xaa3.xa1b.MN0.D xbb1.xa3.M4.D 1.38e-19
C3614 xaa0.xa5.MN2.G xaa0.xa2a.MN0.G 3.32e-19
C3615 xaa6.xe.XA1.MN0.G a_33652_55566# 0.00209f
C3616 AVDD a_34804_54510# 0.00151f
C3617 xaa1.xa4.M0.D m3_37668_116764# 0.074f
C3618 a_5844_60782# li_6204_61812# 1.49e-19
C3619 a_4692_60782# li_4836_61284# 4e-19
C3620 xaa6.xe.XA5.MN0.G a_31132_54158# 1.95e-19
C3621 xaa1.xa3.D m3_4628_70524# 0.0276f
C3622 a_n908_61510# xaa1.xa1.M8.D 0.0251f
C3623 xaa5.xb2_0.MN0.D a_29764_61454# 0.00263f
C3624 AVDD a_n908_61510# 0.00141f
C3625 xaa0.xa5.MN2.G a_n908_55566# 8.96e-19
C3626 a_33652_57326# a_34804_57326# 0.00133f
C3627 xaa6.xf.XA7.MN1.D a_34804_56622# 0.0377f
C3628 xaa6.xc.XA7.MN0.D a_27244_56974# 0.016f
C3629 AVDD a_29764_55566# 0.00151f
C3630 m2_4468_76124# m3_37668_76444# 0.0138f
C3631 xaa3.xa1b.MN0.D li_4836_56708# 0.00345f
C3632 xaa1.xa4.M0.D m1_4468_79004# 67.7f
C3633 a_31132_55566# a_32284_55566# 0.00133f
C3634 xaa6.xd.XA6.MN0.G a_29764_55214# 0.0658f
C3635 xaa6.xd.XA1.MN0.G a_29764_52750# 0.00159f
C3636 xaa6.xe.XA7.MN1.G a_32284_53454# 0.101f
C3637 xaa6.xe.XA7.MP1.G a_31132_53454# 2.78e-19
C3638 a_4692_56206# li_4980_56708# 2e-19
C3639 xaa6.xg.XA7.MN0.D m1_37504_55818# 2.09e-19
C3640 xaa4.xa1.M7.D a_10092_52750# 5.02e-20
C3641 a_36172_53806# a_37324_53806# 0.00133f
C3642 xaa1.xa4.M0.D m3_37748_83164# 0.111f
C3643 li_4468_91484# li_4468_91324# 7.91f
C3644 xaa1.xa3.D a_640_61158# 0.0364f
C3645 xaa5.xa3.xb1_0.G xaa5.xa3.xb1_0.D 0.192f
C3646 xaa5.xb1.MN1.G xaa5.xb2_1.MN0.D 0.0409f
C3647 xaa5.xa3.xb2_0.G a_27244_62510# 0.00184f
C3648 xaa0.xa6.MN0.D xaa1.xa2.M0.D 8.17e-19
C3649 xaa4.xa2.M0.G xaa5.xa4.MN0.D 5.47e-20
C3650 a_356_74698# xaa1.xa3.D 0.00304f
C3651 AVDD a_n908_64150# 0.0038f
C3652 m1_4468_72284# m1_4468_72124# 11.3f
C3653 xaa4.xa2.M0.G xaa4.xa2.M0.D 0.466f
C3654 xaa3.xa1b.MN0.D a_4692_55150# 0.00232f
C3655 a_34804_58030# a_34804_57678# 0.0109f
C3656 PWRUP_1V8 a_29764_56622# 0.0796f
C3657 xaa6.xe.XA1.MN0.G xaa6.xf.XA1.MN0.G 0.0169f
C3658 xaa6.xc.XA1.MN0.G a_28612_57678# 0.0258f
C3659 AVDD a_32284_56622# 0.365f
C3660 a_26092_56270# a_26092_55918# 0.0109f
C3661 xaa6.xe.XA6.MP0.D a_32284_55918# 0.00176f
C3662 xaa6.xd.XA7.MP1.G xaa6.xd.XA3.MP0.D 0.0712f
C3663 xaa6.xf.XA1.MN0.G a_34804_54510# 0.00232f
C3664 xaa6.xc.XA7.MN1.D a_26092_54158# 0.066f
C3665 xaa6.xf.XA7.MP1.G a_34804_54862# 0.029f
C3666 xaa6.xf.XA7.MN1.G a_33652_54862# 0.00608f
C3667 a_31132_56270# xaa6.xe.XA6.MN0.G 0.0677f
C3668 AVDD a_10092_52750# 0.0059f
C3669 xaa1.xa4.M0.D m3_4628_100284# 0.0276f
C3670 a_27244_54510# a_27244_54158# 0.0109f
C3671 xaa6.xg.XA4.MP0.D m1_37504_55818# 0.0264f
C3672 xaa1.xa3.D xaa1.xa2.M8.D 0.0896f
C3673 xaa1.xa4.M0.G a_4692_64126# 0.0799f
C3674 PWRUP_1V8 xaa6.xd.XA7.MN1.D 0.161f
C3675 a_4692_60078# a_5844_60078# 0.00133f
C3676 AVDD xaa6.xe.XA7.MN1.D 1.86f
C3677 xaa4.xa4.M0.D a_10092_55038# 0.0051f
C3678 PWRUP_1V8 a_31132_54510# 0.00467f
C3679 IBPSR_1U xbb1.xa3.M4.D 0.0489f
C3680 xaa1.xa4.M0.D li_4468_112444# 23f
C3681 xaa6.xe.XA1.MN0.G a_32284_55566# 0.0022f
C3682 a_33652_56622# a_34804_56622# 0.00133f
C3683 AVDD a_33652_54510# 0.363f
C3684 xaa6.xf.XA4.MP0.D a_33652_54862# 0.00176f
C3685 a_32284_55214# a_33652_55214# 8.89e-19
C3686 a_26092_55214# a_26092_54862# 0.0109f
C3687 xaa1.xa4.M0.D m3_4788_117564# 0.0138f
C3688 a_5844_60782# li_6132_61812# 4.95e-20
C3689 a_33652_53102# a_33652_52750# 0.0109f
C3690 xbb1.xa3.M4.D a_4308_51918# 1.21e-19
C3691 xaa1.xa3.D m3_37748_70684# 0.111f
C3692 li_4468_75004# li_4468_74204# 39.3f
C3693 li_4468_96284# m1_4468_96284# 23f
C3694 a_26092_61806# a_26092_61454# 0.0109f
C3695 xaa0.xa6.MN0.D xaa0.xa5.MN2.G 0.00284f
C3696 xaa5.xa3.xb1_0.D a_27244_61102# 0.00715f
C3697 xaa5.xb2_0.MN0.D a_28612_61454# 0.00224f
C3698 AVDD a_29764_61806# 0.00139f
C3699 xaa6.xe.XA7.MN1.G xaa6.xe.XA7.MN2.D 0.0148f
C3700 xaa6.xc.XA7.MP1.G a_27244_56974# 0.0291f
C3701 PWRUP_1V8 a_26092_55566# 0.00486f
C3702 xaa0.xa5.MN2.G xaa0.xa1.MN0.G 0.073f
C3703 xaa6.xf.XA7.MN1.D a_33652_56622# 0.0232f
C3704 xaa6.xe.XA1.MN0.G a_34804_56622# 1.73e-19
C3705 xaa6.xc.XA7.MN0.D a_26092_56974# 0.00297f
C3706 AVDD a_28612_55566# 0.383f
C3707 xaa1.xa4.M0.D m1_4468_79964# 67.7f
C3708 xaa6.xd.XA6.MN0.G a_28612_55214# 0.0827f
C3709 xaa6.xd.XA7.MN1.D a_29764_52750# 6.12e-22
C3710 xaa6.xe.XA7.MN1.G a_31132_53454# 0.015f
C3711 a_4692_56206# li_4836_56708# 4e-19
C3712 a_5844_56206# li_6204_57236# 1.49e-19
C3713 xaa6.xg.XA7.MP1.G m1_37504_55818# 0.242f
C3714 xaa6.xg.XA7.MN0.D m1_37504_57930# 0.0293f
C3715 a_29764_53806# xaa6.xd.XA1.MN0.D 0.00176f
C3716 xaa1.xa4.M0.D m3_37668_83164# 0.074f
C3717 xaa5.xa3.xb2_0.G a_26092_62510# 0.00665f
C3718 xaa4.xa2.M0.G a_29764_62510# 3.48e-19
C3719 xaa5.xb2_4.MN0.D CK 7.29e-20
C3720 xaa3.xa5a.MN0.D a_5844_62366# 0.0766f
C3721 IBPSR_1U xaa1.xa2.M2.D 0.026f
C3722 AVDD a_29764_64270# 0.00139f
C3723 m1_4468_99164# m2_4468_99164# 12.9f
C3724 IBPSR_1U a_4692_55150# 0.00178f
C3725 xaa3.xa1b.MN0.D a_5844_55502# 0.00224f
C3726 a_27244_58030# xaa6.xc.XA7.MP1.G 3.8e-19
C3727 PWRUP_1V8 a_28612_56622# 0.0658f
C3728 xaa6.xc.XA1.MN0.G a_27244_57678# 0.00249f
C3729 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN1.D 0.274f
C3730 AVDD a_31132_56622# 0.00151f
C3731 a_4692_55854# a_4692_55502# 0.0109f
C3732 xaa6.xf.XA1.MN0.G a_33652_54510# 1.17e-19
C3733 xaa6.xf.XA7.MN1.D a_34804_54510# 0.072f
C3734 xaa1.xa4.M0.D li_4468_78844# 23f
C3735 xaa6.xf.XA7.MP1.G a_33652_54862# 0.0986f
C3736 xaa6.xf.XA7.MN1.G a_32284_54862# 7.1e-20
C3737 a_34804_56270# a_36172_56270# 8.89e-19
C3738 xaa1.xa4.M0.D m3_37748_100444# 0.111f
C3739 a_34804_54510# a_36172_54510# 8.89e-19
C3740 xaa6.xf.XA3.MP0.D a_33652_54158# 0.00176f
C3741 li_4468_108764# li_4468_108604# 7.91f
C3742 PWRUP_1V8 xaa6.xc.XA1.MN0.G 0.212f
C3743 AVDD xaa6.xd.XA1.MN0.G 1.64f
C3744 PWRUP_1V8 a_29764_54510# 0.00467f
C3745 IBPSR_1U xaa4.xa1.M0.D 0.0279f
C3746 xaa0.xa5.MN2.G a_n908_54862# 2.88e-19
C3747 xaa6.xe.XA7.MN1.D a_32284_55566# 0.00147f
C3748 xaa6.xg.XA7.MN0.D xaa6.xg.XA6.MN0.G 1.04e-19
C3749 a_28612_57326# xaa6.xd.XA6.MN0.G 5e-20
C3750 xaa6.xe.XA1.MN0.G a_31132_55566# 1.25e-19
C3751 xaa6.xe.XA7.MN1.G a_33652_55918# 7.1e-20
C3752 xaa6.xe.XA7.MP1.G a_32284_55918# 0.0292f
C3753 AVDD a_32284_54510# 0.363f
C3754 xaa1.xa4.M0.D m3_4628_117564# 0.0276f
C3755 xaa6.xd.XA5.MN0.G a_29764_54158# 1.95e-19
C3756 xaa6.xg.XA6.MP0.D m1_37504_55818# 0.00192f
C3757 xaa1.xa3.D m3_37668_70684# 0.074f
C3758 a_n908_61510# a_640_61510# 6.96e-19
C3759 a_29764_61806# xaa5.xb1.MN1.D 0.0682f
C3760 xaa5.xa3.xb1_0.D a_26092_61102# 0.0561f
C3761 xaa3.xa5a.MN0.D a_5844_60078# 7.03e-19
C3762 AVDD a_28612_61806# 0.352f
C3763 m2_4468_117404# m3_37748_117724# 0.0138f
C3764 a_32284_57326# a_33652_57326# 8.89e-19
C3765 xaa6.xc.XA7.MP1.G a_26092_56974# 2.35e-19
C3766 xaa6.xc.XA7.MN1.G a_27244_56974# 0.0035f
C3767 xaa0.xa5.MN2.G a_244_55918# 0.0674f
C3768 xaa6.xe.XA1.MN0.G a_33652_56622# 0.00369f
C3769 AVDD a_27244_55566# 0.383f
C3770 xaa6.xg.XA7.MN1.D a_37324_53102# 5.24e-20
C3771 xaa1.xa4.M0.D m1_4468_80924# 67.7f
C3772 xaa6.xg.XA5.MN0.G a_37324_55566# 0.0889f
C3773 a_29764_55566# a_31132_55566# 8.89e-19
C3774 xaa6.xg.XA7.MN1.G xaa6.xg.XA1.MN0.D 7.79e-19
C3775 xaa6.xd.XA7.MN1.D a_28612_52750# 3.67e-21
C3776 a_5844_56206# li_6132_57236# 4.95e-20
C3777 xaa6.xg.XA7.MN1.G m1_37504_55818# 0.153f
C3778 xaa6.xg.XA7.MP1.G m1_37504_57930# 0.13f
C3779 a_34804_53806# a_36172_53806# 8.89e-19
C3780 xaa6.xg.XA3.MN1.G a_37324_52750# 1.28e-19
C3781 xaa1.xa4.M0.D m3_4788_83964# 0.0138f
C3782 li_4468_92284# li_4468_91484# 39.3f
C3783 xaa4.xa2.M0.G a_28612_62510# 0.0362f
C3784 xaa5.xa3.xb2_0.G xaa5.xb2_2.MN0.D 0.00451f
C3785 a_29764_63566# CK 3.97e-20
C3786 xaa3.xa5a.MN0.D a_4692_62366# 0.0913f
C3787 xaa5.xb2_4.MN0.D a_29764_62862# 0.00263f
C3788 a_n908_63270# xaa1.xa2.M2.D 8.62e-20
C3789 AVDD a_28612_64270# 0.351f
C3790 xaa3.xa1b.MN0.D a_4692_55502# 0.00861f
C3791 xaa6.xc.XA7.MN1.D a_27244_57678# 0.0893f
C3792 a_33652_58030# a_33652_57678# 0.0109f
C3793 xaa0.xa5.MN2.G a_28612_57678# 2.93e-19
C3794 a_27244_58030# xaa6.xc.XA7.MN1.G 3.89e-19
C3795 PWRUP_1V8 a_27244_56622# 0.0674f
C3796 xaa6.xe.XA7.MN1.D xaa6.xf.XA7.MN1.D 0.00435f
C3797 xaa6.xc.XA1.MN0.G a_26092_57678# 1.35e-19
C3798 AVDD a_29764_56622# 0.00151f
C3799 xaa6.xe.XA6.MN0.D a_31132_55918# 0.00176f
C3800 PWRUP_1V8 a_34804_53102# 1.28e-19
C3801 a_29764_56270# xaa6.xd.XA6.MN0.G 0.0661f
C3802 xaa6.xf.XA7.MN1.D a_33652_54510# 0.0851f
C3803 xaa6.xe.XA1.MN0.G a_34804_54510# 1.02e-19
C3804 AVDD a_37324_53102# 0.485f
C3805 xaa1.xa4.M0.D m3_37668_100444# 0.074f
C3806 a_26092_54510# a_26092_54158# 0.0109f
C3807 xaa4.xa2.M0.G m3_22620_52900# 0.0273f
C3808 xaa6.xg.XA4.MP1.G m1_37504_55818# 0.0171f
C3809 a_n908_64150# xaa1.xa4.M0.G 0.073f
C3810 li_4468_74204# m1_4468_74204# 23f
C3811 PWRUP_1V8 xaa6.xc.XA7.MN1.D 0.162f
C3812 xaa1.xa1.M2.D a_n908_59750# 2.99e-19
C3813 xaa3.xa3a.MN0.D a_5844_60078# 0.0766f
C3814 AVDD xaa6.xd.XA7.MN1.D 1.86f
C3815 m2_4468_103964# m3_37748_104284# 0.0138f
C3816 xaa6.xg.XA7.MP1.G xaa6.xg.XA6.MN0.G 0.111f
C3817 xaa1.xa4.M0.D li_4468_113404# 23f
C3818 xaa6.xe.XA7.MN1.D a_31132_55566# 0.00699f
C3819 a_32284_56622# a_33652_56622# 8.89e-19
C3820 xaa6.xd.XA1.MN0.G a_32284_55566# 1.11e-19
C3821 xaa6.xe.XA7.MN1.G a_32284_55918# 0.00733f
C3822 xaa6.xe.XA7.MP1.G a_31132_55918# 0.0294f
C3823 AVDD a_31132_54510# 0.00151f
C3824 xaa6.xe.XA4.MP0.D a_32284_54862# 0.00176f
C3825 a_31132_55214# a_32284_55214# 0.00133f
C3826 xaa1.xa4.M0.D m3_37748_117724# 0.111f
C3827 xaa6.xd.XA5.MN0.G a_28612_54158# 1.28e-19
C3828 a_32284_53102# a_32284_52750# 0.0109f
C3829 a_10092_52750# a_11712_52750# 6.4e-19
C3830 xaa6.xg.XA6.MP0.D m1_37504_57930# 4.24e-20
C3831 xaa1.xa3.D m3_4788_71484# 0.0138f
C3832 li_4468_75164# li_4468_75004# 7.91f
C3833 xaa1.xa2.M0.D PWRUP_1V8 0.00408f
C3834 xaa5.xa3.xc2a.D a_27244_61454# 0.00176f
C3835 a_28612_61806# xaa5.xb1.MN1.D 0.0674f
C3836 xaa3.xa5a.MN0.D a_4692_60078# 1.15e-19
C3837 AVDD a_27244_61806# 0.364f
C3838 m2_4468_117404# m3_37668_117724# 0.0138f
C3839 xaa6.xc.XA7.MN1.G a_26092_56974# 0.00922f
C3840 xaa4.xa2.M0.G a_10092_54510# 0.0705f
C3841 PWRUP_1V8 xaa6.xg.XA5.MN0.G 0.0749f
C3842 xaa0.xa5.MN2.G a_n908_55918# 0.0659f
C3843 xaa6.xe.XA1.MN0.G a_32284_56622# 0.0022f
C3844 xaa6.xd.XA7.MN0.D xaa6.xd.XA7.MN2.D 0.0618f
C3845 AVDD a_26092_55566# 0.00159f
C3846 xaa6.xg.XA7.MN1.D a_36172_53102# 8.73e-21
C3847 xaa3.xa1b.MN0.D li_4980_58996# 2.55e-19
C3848 xaa1.xa4.M0.D m1_4468_81884# 67.7f
C3849 xaa6.xg.XA5.MN0.G a_36172_55566# 0.112f
C3850 xaa6.xc.XA6.MN0.G a_27244_55214# 0.0811f
C3851 xaa6.xg.XA5.MN0.D a_37324_55566# 0.00224f
C3852 xaa6.xg.XA7.MN1.G m1_37504_57930# 0.00933f
C3853 a_4308_53678# xbb1.xa3.M5.D 2.99e-19
C3854 xaa6.xg.XA3.MN1.G a_36172_52750# 2.64e-19
C3855 xaa1.xa4.M0.D m3_4628_83964# 0.0276f
C3856 AVDD xaa5.xb3.MP1.D 0.476f
C3857 xaa5.xa3.xb2_0.G xaa5.xa3.xb2_0.D 0.145f
C3858 xaa5.xb1.MN1.G a_29764_62510# 0.00547f
C3859 xaa0.xa6.MN0.D xaa1.xa2.M1.D 8.17e-19
C3860 xaa4.xa2.M0.G a_27244_62510# 6.38e-19
C3861 a_5844_62718# a_5844_62366# 0.0109f
C3862 xaa5.xb2_4.MN0.D a_28612_62862# 0.00224f
C3863 m1_4468_100124# m2_4468_100124# 12.9f
C3864 xaa6.xd.XA1.MN0.G xaa6.xf.XA7.MN1.D 4.33e-19
C3865 IBPSR_1U a_4692_55502# 7.97e-19
C3866 xaa0.xa5.MN2.G a_27244_57678# 0.0209f
C3867 xaa6.xc.XA7.MN1.D a_26092_57678# 0.132f
C3868 a_26092_58030# xaa6.xc.XA7.MN1.G 0.00215f
C3869 PWRUP_1V8 a_26092_56622# 0.0777f
C3870 xaa6.xe.XA7.MN1.D xaa6.xe.XA1.MN0.G 0.0209f
C3871 AVDD a_28612_56622# 0.365f
C3872 m2_4468_90524# m3_37748_90844# 0.0138f
C3873 xaa1.xa4.M0.D li_4468_79804# 23f
C3874 xaa6.xc.XA7.MP1.G xaa6.xc.XA3.MP0.D 0.0712f
C3875 a_33652_56270# a_34804_56270# 0.00133f
C3876 a_28612_56270# xaa6.xd.XA6.MN0.G 0.0735f
C3877 xaa6.xg.XA6.MP0.D xaa6.xg.XA6.MN0.G 0.0093f
C3878 xaa6.xe.XA1.MN0.G a_33652_54510# 0.00196f
C3879 AVDD a_36172_53102# 0.00163f
C3880 xaa1.xa4.M0.D m3_4788_101244# 0.0138f
C3881 a_33652_54510# a_34804_54510# 0.00133f
C3882 xaa6.xe.XA3.MP0.D a_32284_54158# 0.00176f
C3883 xaa4.xa2.M0.G m3_22548_52900# 0.0137f
C3884 li_4468_109564# li_4468_108764# 39.3f
C3885 xaa1.xa3.D xaa0.xa6.MN0.D 0.0217f
C3886 PWRUP_1V8 xaa0.xa5.MN2.G 5.41f
C3887 xaa3.xa3a.MN0.D a_4692_60078# 0.0913f
C3888 AVDD xaa6.xc.XA1.MN0.G 3.51f
C3889 m2_4468_103964# m3_37668_104284# 0.0138f
C3890 xaa6.xg.XA7.MN1.G xaa6.xg.XA6.MN0.G 0.0417f
C3891 a_27244_57326# xaa6.xc.XA6.MN0.G 5e-20
C3892 xaa6.xd.XA1.MN0.G a_31132_55566# 0.00205f
C3893 xaa6.xe.XA7.MN1.G a_31132_55918# 7.37e-19
C3894 AVDD a_29764_54510# 0.00151f
C3895 xaa4.xa1.M8.D xaa4.xa1.M7.D 0.0488f
C3896 xaa6.xg.XA4.MP0.D xaa6.xg.XA4.MN0.G 0.0093f
C3897 xaa1.xa4.M0.D m3_37668_117724# 0.074f
C3898 xaa1.xa3.D m3_4628_71484# 0.0276f
C3899 li_4468_97244# m1_4468_97244# 23f
C3900 xaa5.xb2_0.MN0.D PWRUP_1V8 5.71e-20
C3901 AVDD a_26092_61806# 0.00159f
C3902 PWRUP_1V8 xaa6.xg.XA5.MN0.D 0.00139f
C3903 a_31132_57326# a_32284_57326# 0.00133f
C3904 xaa3.xa1capd.B a_5844_55854# 0.00414f
C3905 a_5844_57790# a_5844_56206# 0.00744f
C3906 xaa0.xa5.MN2.G xaa0.xa5.MP1.D 0.00991f
C3907 xaa6.xe.XA7.MN1.D a_32284_56622# 0.0232f
C3908 xaa6.xe.XA1.MN0.G a_31132_56622# 1.25e-19
C3909 xaa6.xd.XA7.MN1.G xaa6.xd.XA7.MN2.D 0.0148f
C3910 AVDD xaa4.xa1.M8.D 0.077f
C3911 m2_4468_77084# m3_37748_77404# 0.0138f
C3912 xaa3.xa1b.MN0.D li_4836_58996# 0.00265f
C3913 xaa1.xa4.M0.D m1_4468_82844# 67.7f
C3914 xaa6.xd.XA7.MN1.G a_29764_53454# 0.015f
C3915 xaa6.xc.XA6.MN0.G a_26092_55214# 0.0674f
C3916 xaa6.xg.XA5.MN0.D a_36172_55566# 0.00224f
C3917 xaa6.xc.XA1.MN0.G a_27244_52750# 0.00177f
C3918 a_28612_55566# a_29764_55566# 0.00133f
C3919 a_33652_53806# a_34804_53806# 0.00133f
C3920 xaa1.xa4.M0.D m3_37748_84124# 0.111f
C3921 li_4468_92444# li_4468_92284# 7.91f
C3922 xaa1.xa2.M4.D xaa1.xa2.M3.D 0.0488f
C3923 xaa5.xb1.MN1.G a_28612_62510# 9.6e-19
C3924 xaa5.xa3.xb2_0.G CK 0.0589f
C3925 AVDD a_29764_64622# 0.00584f
C3926 a_n508_74698# xaa1.xa3.D 0.00272f
C3927 xaa6.xd.XA1.MN0.G xaa6.xe.XA1.MN0.G 0.071f
C3928 IBPSR_1U xaa4.xa2.M0.D 0.0205f
C3929 xaa0.xa5.MN2.G a_26092_57678# 0.00456f
C3930 a_32284_58030# a_32284_57678# 0.0109f
C3931 PWRUP_1V8 a_37324_56974# 0.0658f
C3932 AVDD a_27244_56622# 0.365f
C3933 m2_4468_90524# m3_37668_90844# 0.0138f
C3934 xaa6.xe.XA7.MP1.G a_32284_54862# 0.097f
C3935 xaa6.xe.XA7.MN1.G a_33652_54862# 7.1e-20
C3936 xaa6.xd.XA6.MN0.D a_29764_55918# 0.00176f
C3937 xaa4.xa4.M0.D xaa4.xa1.M3.D 4.85e-19
C3938 xaa6.xc.XA7.MP1.G xaa6.xc.XA3.MN0.D 0.0472f
C3939 xaa6.xc.XA7.MN1.G xaa6.xc.XA3.MP0.D 0.00252f
C3940 xaa6.xg.XA6.MN0.D xaa6.xg.XA6.MN0.G 0.0093f
C3941 xaa6.xe.XA1.MN0.G a_32284_54510# 0.00267f
C3942 xaa6.xg.XA7.MP1.G xaa6.xg.XA4.MN0.G 0.127f
C3943 AVDD a_34804_53102# 0.00163f
C3944 xaa1.xa4.M0.D m3_4628_101244# 0.0276f
C3945 xaa4.xa2.M0.G m3_13116_53076# 0.0634f
C3946 xaa1.xa3.D a_n908_63622# 0.0276f
C3947 PWRUP_1V8 a_37324_58030# 8.58e-19
C3948 AVDD xaa6.xc.XA7.MN1.D 1.86f
C3949 xaa6.xg.XA7.MN1.D xaa6.xg.XA5.MN0.G 0.29f
C3950 PWRUP_1V8 a_26092_54510# 0.0046f
C3951 xaa1.xa4.M0.D li_4468_114364# 23f
C3952 a_31132_56622# a_32284_56622# 0.00133f
C3953 xaa6.xd.XA1.MN0.G a_29764_55566# 0.00217f
C3954 AVDD a_28612_54510# 0.363f
C3955 xaa6.xe.XA4.MN0.D a_31132_54862# 0.00176f
C3956 xaa6.xg.XA4.MP0.D a_37324_55214# 0.0467f
C3957 a_29764_55214# a_31132_55214# 8.89e-19
C3958 xaa6.xg.XA4.MN0.D xaa6.xg.XA4.MN0.G 0.0093f
C3959 xaa6.xc.XA5.MN0.G a_27244_54158# 1.28e-19
C3960 xaa1.xa3.D m3_37748_71644# 0.111f
C3961 a_31132_53102# a_31132_52750# 0.0109f
C3962 li_4468_75964# li_4468_75164# 39.3f
C3963 xaa1.xa2.M0.D xaa1.xa1.M8.D 0.00584f
C3964 xaa3.xa1b.MN0.D a_4692_57790# 0.00455f
C3965 xaa3.xa5a.MN0.D xaa3.xa3a.MN0.D 0.00369f
C3966 PWRUP_1V8 xaa6.xf.XA5.MN0.G 0.0755f
C3967 xaa6.xg.XA7.MN0.D a_37324_57326# 0.0525f
C3968 xaa6.xd.XA1.MN0.G a_32284_56622# 0.00119f
C3969 xaa3.xa1capd.B a_4692_55854# 0.00429f
C3970 xaa6.xe.XA7.MN1.D a_31132_56622# 0.0377f
C3971 AVDD xaa6.xg.XA5.MN0.G 0.879f
C3972 m2_4468_77084# m3_37668_77404# 0.0138f
C3973 xaa6.xf.XA7.MN1.G xaa6.xf.XA1.MN0.D 0.123f
C3974 xaa6.xc.XA7.MN1.D a_27244_52750# 3.67e-21
C3975 xaa6.xf.XA1.MN0.G a_34804_53102# 0.0721f
C3976 xaa6.xd.XA7.MN1.G a_28612_53454# 0.101f
C3977 xaa6.xd.XA7.MP1.G a_29764_53454# 2.78e-19
C3978 xaa6.xc.XA1.MN0.G a_26092_52750# 0.00263f
C3979 xaa1.xa4.M0.D m1_4468_83804# 67.7f
C3980 a_26092_53806# xaa6.xc.XA1.MN0.D 0.00176f
C3981 xaa1.xa4.M0.D m3_37668_84124# 0.074f
C3982 a_4692_62718# a_4692_62366# 0.0109f
C3983 xaa5.xa3.xb1_0.G a_26092_62510# 0.00235f
C3984 xaa4.xa2.M0.G xaa5.xb2_2.MN0.D 0.174f
C3985 a_29764_63918# CK 3.54e-19
C3986 xaa5.xa3.xb2_0.G a_29764_62862# 3.89e-19
C3987 AVDD a_28612_64622# 0.335f
C3988 m1_4468_101084# m2_4468_101084# 12.9f
C3989 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN1.D 0.262f
C3990 AVDD a_26092_56622# 0.00159f
C3991 PWRUP_1V8 a_36172_56974# 0.0768f
C3992 a_36172_56622# xaa6.xg.XA5.MN0.G 6.14e-19
C3993 xaa6.xe.XA7.MP1.G a_31132_54862# 0.029f
C3994 xaa6.xe.XA7.MN1.G a_32284_54862# 0.00608f
C3995 xaa1.xa4.M0.D li_4468_80764# 23f
C3996 xaa4.xa4.M0.D xaa4.xa1.M4.D 5.29e-19
C3997 xaa6.xc.XA7.MN1.G xaa6.xc.XA3.MN0.D 0.0288f
C3998 a_32284_56270# a_33652_56270# 8.89e-19
C3999 a_27244_56270# xaa6.xc.XA6.MN0.G 0.0719f
C4000 xaa6.xe.XA7.MN1.D a_32284_54510# 0.0836f
C4001 xaa6.xe.XA1.MN0.G a_31132_54510# 6.72e-19
C4002 xaa6.xg.XA7.MN1.G xaa6.xg.XA4.MN0.G 0.014f
C4003 xaa6.xg.XA7.MP1.G a_37324_55214# 0.027f
C4004 AVDD a_33652_53102# 0.488f
C4005 xaa6.xe.XA3.MN0.D a_31132_54158# 0.00176f
C4006 a_32284_54510# a_33652_54510# 8.89e-19
C4007 xaa1.xa4.M0.D m3_37748_101404# 0.111f
C4008 xaa4.xa2.M0.G m3_13044_53076# 0.106f
C4009 li_4468_109724# li_4468_109564# 7.91f
C4010 li_4468_75164# m1_4468_75164# 23f
C4011 PWRUP_1V8 a_36172_58030# 0.00223f
C4012 AVDD xaa0.xa5.MN2.G 3.37f
C4013 xaa6.xf.XA1.MN0.G xaa6.xg.XA5.MN0.G 0.00846f
C4014 a_37324_56974# a_37324_56622# 0.0109f
C4015 xaa6.xd.XA7.MN1.D a_29764_55566# 0.00699f
C4016 xaa6.xf.XA7.MN0.D xaa6.xf.XA6.MN0.G 3.13e-19
C4017 xaa6.xd.XA1.MN0.G a_28612_55566# 1.35e-19
C4018 xaa6.xg.XA7.MN1.D xaa6.xg.XA5.MN0.D 0.0864f
C4019 AVDD a_27244_54510# 0.363f
C4020 xaa6.xg.XA5.MN0.G a_37324_54510# 0.00224f
C4021 xaa6.xg.XA4.MP1.G xaa6.xg.XA4.MN0.G 0.0184f
C4022 xaa6.xc.XA5.MN0.G a_26092_54158# 1.95e-19
C4023 xaa1.xa3.D m3_37668_71644# 0.074f
C4024 xaa1.xa2.M1.D PWRUP_1V8 0.00279f
C4025 a_28612_61806# a_29764_61806# 0.00133f
C4026 IBPSR_1U a_4692_57790# 1.59e-20
C4027 xaa3.xa1b.MN0.D xaa3.xa1capd.B 0.406f
C4028 xaa5.xa3.xb1_0.D xaa5.xa3.xc1a.D 0.0802f
C4029 AVDD xaa5.xb2_0.MN0.D 0.55f
C4030 a_29764_57326# a_31132_57326# 8.89e-19
C4031 xaa6.xg.XA7.MN0.D a_36172_57326# 0.055f
C4032 xaa6.xd.XA1.MN0.G a_31132_56622# 0.00133f
C4033 xaa6.xg.XA7.MN1.D a_37324_56974# 0.00166f
C4034 xaa3.xa1capd.B a_5844_56206# 0.0536f
C4035 a_4692_57790# a_4692_56206# 0.00744f
C4036 xaa6.xg.XA7.MP1.G a_37324_57326# 0.0964f
C4037 PWRUP_1V8 xaa6.xe.XA5.MN0.G 0.0749f
C4038 AVDD xaa6.xg.XA5.MN0.D 0.216f
C4039 xaa6.xc.XA7.MN1.D a_26092_52750# 6.12e-22
C4040 xaa6.xf.XA1.MN0.G a_33652_53102# 0.0658f
C4041 xaa6.xf.XA7.MN1.D a_34804_53102# 8.73e-21
C4042 xaa6.xd.XA7.MN1.G a_27244_53454# 7.1e-20
C4043 xaa6.xd.XA7.MP1.G a_28612_53454# 1.07e-19
C4044 xaa6.xf.XA6.MN0.G xaa6.xf.XA4.MN0.D 0.0093f
C4045 xaa6.xf.XA5.MN0.G a_34804_55566# 0.113f
C4046 a_27244_55566# a_28612_55566# 8.89e-19
C4047 xaa1.xa4.M0.D m1_4468_84764# 67.7f
C4048 a_32284_53806# a_33652_53806# 8.89e-19
C4049 xaa1.xa4.M0.D m3_4788_84924# 0.0138f
C4050 li_4468_93244# li_4468_92444# 39.3f
C4051 xaa3.xa6.MN0.D a_5844_62366# 0.00224f
C4052 a_5844_62718# xaa3.xa5a.MN0.D 0.0658f
C4053 xaa5.xb2_4.MN0.D xaa5.xb2_3.MN0.D 0.197f
C4054 xaa1.xa3.D PWRUP_1V8 0.0281f
C4055 a_28612_63918# CK 4.49e-19
C4056 xaa5.xa3.xb2_0.G a_28612_62862# 0.00172f
C4057 xaa4.xa2.M0.G xaa5.xa3.xb2_0.D 0.0044f
C4058 xbb0.xa1.XA1.N xaa1.xa3.D 0.0687f
C4059 xaa6.xd.XA7.MN1.D xaa6.xe.XA7.MN1.D 0.00642f
C4060 a_37324_58030# xaa6.xg.XA7.MN1.D 0.0658f
C4061 a_31132_58030# a_31132_57678# 0.0109f
C4062 AVDD a_37324_56974# 0.405f
C4063 PWRUP_1V8 a_34804_56974# 0.0755f
C4064 xaa6.xe.XA7.MN1.G a_31132_54862# 0.0724f
C4065 xaa6.xd.XA1.MN0.G a_32284_54510# 1.11e-19
C4066 xaa6.xd.XA6.MP0.D a_28612_55918# 0.00176f
C4067 PWRUP_1V8 a_29764_53102# 1.28e-19
C4068 a_26092_56270# xaa6.xc.XA6.MN0.G 0.0677f
C4069 xaa6.xf.XA6.MN0.D xaa6.xf.XA6.MN0.G 0.0093f
C4070 xaa6.xe.XA7.MN1.D a_31132_54510# 0.0736f
C4071 xaa6.xg.XA7.MN1.G a_37324_55214# 0.00688f
C4072 xaa6.xg.XA7.MP1.G a_36172_55214# 0.0944f
C4073 AVDD a_32284_53102# 0.486f
C4074 xaa1.xa4.M0.D m3_37668_101404# 0.074f
C4075 xaa4.xa2.M0.G m3_22620_53956# 0.0273f
C4076 a_28612_64270# a_29764_64270# 0.00133f
C4077 xaa1.xa1.M3.D a_n908_59750# 1.81e-19
C4078 a_640_60278# xaa1.xb1.M0.D 0.00155f
C4079 a_5844_60430# a_5844_60078# 0.0109f
C4080 PWRUP_1V8 a_34804_58030# 0.00639f
C4081 AVDD a_37324_58030# 0.344f
C4082 xaa6.xf.XA1.MN0.G xaa6.xg.XA5.MN0.D 0.00222f
C4083 xaa6.xd.XA7.MN1.G a_29764_55918# 7.37e-19
C4084 a_29764_56622# a_31132_56622# 8.89e-19
C4085 xaa6.xd.XA7.MN1.D a_28612_55566# 0.00147f
C4086 xaa6.xf.XA7.MN1.G xaa6.xf.XA6.MN0.G 0.329f
C4087 xaa6.xc.XA1.MN0.G a_29764_55566# 1.02e-19
C4088 AVDD a_26092_54510# 0.00159f
C4089 xaa1.xa4.M0.D li_4468_115324# 23f
C4090 xaa6.xg.XA5.MN0.G a_36172_54510# 0.00236f
C4091 xaa6.xd.XA4.MN0.D a_29764_54862# 0.00176f
C4092 xaa6.xg.XA4.MN0.D a_36172_55214# 0.0472f
C4093 a_28612_55214# a_29764_55214# 0.00133f
C4094 xaa6.xg.XA4.MP1.G a_37324_55214# 0.0674f
C4095 a_29764_53102# a_29764_52750# 0.0109f
C4096 li_4468_76124# li_4468_75964# 7.91f
C4097 li_4468_98204# m1_4468_98204# 23f
C4098 a_29764_62158# PWRUP_1V8 2.56e-20
C4099 xaa5.xb2_0.MN0.D xaa5.xb1.MN1.D 0.184f
C4100 IBPSR_1U xaa3.xa1capd.B 3.88e-20
C4101 CK a_29764_61102# 3.97e-20
C4102 AVDD xaa5.xa3.xc2a.D 0.159f
C4103 m1_4468_69404# m2_4468_69404# 12.9f
C4104 xaa6.xd.XA1.MN0.G a_29764_56622# 0.00134f
C4105 xaa6.xg.XA7.MN1.D a_36172_56974# 0.0092f
C4106 IBPSR_1U a_10092_54510# 0.0677f
C4107 xaa3.xa1capd.B a_4692_56206# 0.0583f
C4108 xaa6.xc.XA7.MN0.D xaa6.xc.XA7.MN2.D 0.0618f
C4109 xaa6.xg.XA7.MP1.G a_36172_57326# 9.02e-20
C4110 xaa6.xg.XA7.MN1.G a_37324_57326# 0.00186f
C4111 PWRUP_1V8 xaa6.xd.XA5.MN0.G 0.0755f
C4112 AVDD xaa6.xf.XA5.MN0.G 0.88f
C4113 xaa3.xa1b.MN0.D li_4980_61284# 2.55e-19
C4114 xaa6.xf.XA7.MN1.D a_33652_53102# 5.24e-20
C4115 xaa6.xf.XA6.MN0.G xaa6.xf.XA4.MP0.D 0.0357f
C4116 xaa6.xf.XA5.MN0.G a_33652_55566# 0.0873f
C4117 xaa1.xa4.M0.D m1_4468_85724# 67.7f
C4118 xbb1.xa3.M7.D xbb1.xa3.M6.D 0.0488f
C4119 xaa1.xa4.M0.D m3_4628_84924# 0.0276f
C4120 xaa3.xa6.MN0.D a_4692_62366# 0.00346f
C4121 a_4692_62718# xaa3.xa5a.MN0.D 0.0728f
C4122 xaa5.xb2_4.MN0.D a_29764_63214# 0.126f
C4123 xaa5.xb1.MN1.G xaa5.xb2_2.MN0.D 0.0405f
C4124 xaa5.xa3.xb1_0.G xaa5.xa3.xb2_0.D 0.0181f
C4125 xaa4.xa2.M0.G CK 0.794f
C4126 xaa5.xa3.xb2_0.G a_27244_62862# 0.00266f
C4127 a_n940_74698# xaa1.xa3.D 0.00106f
C4128 m1_4468_102044# m2_4468_102044# 12.9f
C4129 xaa6.xc.XA1.MN0.G xaa6.xe.XA7.MN1.D 2.06e-19
C4130 xaa6.xd.XA7.MN1.D xaa6.xd.XA1.MN0.G 0.0169f
C4131 a_36172_58030# xaa6.xg.XA7.MN1.D 0.0711f
C4132 a_37324_58030# xaa6.xf.XA1.MN0.G 0.0227f
C4133 PWRUP_1V8 a_33652_56974# 0.0674f
C4134 AVDD a_36172_56974# 0.00151f
C4135 xaa6.xd.XA1.MN0.G a_31132_54510# 0.00193f
C4136 xaa1.xa4.M0.D li_4468_81724# 23f
C4137 xaa6.xg.XA7.MN1.D xaa6.xg.XA3.MP0.D 0.0844f
C4138 a_31132_56270# a_32284_56270# 0.00133f
C4139 xaa6.xf.XA6.MP0.D xaa6.xf.XA6.MN0.G 0.0116f
C4140 xaa6.xg.XA7.MN1.G a_36172_55214# 1.97e-19
C4141 AVDD a_31132_53102# 0.00163f
C4142 xaa6.xd.XA3.MN0.D a_29764_54158# 0.00176f
C4143 a_31132_54510# a_32284_54510# 0.00133f
C4144 xaa1.xa4.M0.D m3_4788_102204# 0.0138f
C4145 xaa4.xa2.M0.G m3_22548_53956# 0.0137f
C4146 li_4468_110524# li_4468_109724# 39.3f
C4147 PWRUP_1V8 a_33652_58030# 4.25e-19
C4148 AVDD a_36172_58030# 0.00519f
C4149 m2_4468_104924# m3_37748_105244# 0.0138f
C4150 xaa6.xg.XA7.MP1.G a_37324_56270# 0.0268f
C4151 xaa6.xf.XA1.MN0.G xaa6.xf.XA5.MN0.G 0.00917f
C4152 PWRUP_1V8 xaa6.xg.XA3.MN1.G 0.382f
C4153 xaa6.xd.XA7.MP1.G a_29764_55918# 0.0294f
C4154 xaa6.xd.XA7.MN1.G a_28612_55918# 0.00733f
C4155 a_36172_56974# a_36172_56622# 0.0109f
C4156 xaa6.xc.XA1.MN0.G a_28612_55566# 0.00209f
C4157 xaa6.xf.XA7.MP1.G xaa6.xf.XA6.MN0.G 0.524f
C4158 xaa6.xf.XA7.MN1.G xaa6.xe.XA6.MN0.G 3.47e-19
C4159 AVDD xaa6.xg.XA3.MP0.D 0.133f
C4160 a_36172_55566# xaa6.xg.XA3.MN1.G 4.21e-19
C4161 a_2948_74698# m2_4468_74204# 7.48e-19
C4162 xaa1.xa4.M0.D m2_4468_72284# 59.5f
C4163 xaa1.xa2.M1.D xaa1.xa1.M8.D 0.00304f
C4164 xaa1.xa2.M0.D a_n908_61510# 0.00155f
C4165 a_27244_61806# a_28612_61806# 8.89e-19
C4166 xaa3.xa1b.MN0.D a_4692_58142# 0.00455f
C4167 xaa5.xa3.xb2_0.D a_27244_61102# 0.164f
C4168 a_28612_57326# a_29764_57326# 0.00133f
C4169 xaa6.xd.XA7.MN1.D a_29764_56622# 0.0377f
C4170 xaa6.xg.XA7.MN1.D a_34804_56974# 1.31e-19
C4171 xaa6.xf.XA1.MN0.G a_36172_56974# 0.00138f
C4172 xaa6.xg.XA7.MN1.G a_36172_57326# 0.0781f
C4173 PWRUP_1V8 xaa6.xc.XA5.MN0.G 0.0747f
C4174 AVDD xaa6.xe.XA5.MN0.G 0.88f
C4175 xaa0.xa5.MN2.G a_11712_52750# 3.98e-19
C4176 xaa6.xg.XA7.MP1.G a_37324_53806# 0.00282f
C4177 a_26092_55566# a_27244_55566# 0.00133f
C4178 xaa1.xa4.M0.D m1_4468_86684# 67.7f
C4179 xaa3.xa1b.MN0.D li_4836_61284# 0.00265f
C4180 a_31132_53806# a_32284_53806# 0.00133f
C4181 xaa1.xa4.M0.D m3_37748_85084# 0.111f
C4182 li_4468_93404# li_4468_93244# 7.91f
C4183 xaa5.xb2_4.MN0.D a_28612_63214# 0.0878f
C4184 a_29764_63566# a_29764_63214# 0.0109f
C4185 xaa0.xa6.MN0.D xaa1.xa2.M2.D 8.17e-19
C4186 xaa1.xa3.D xaa1.xa1.M8.D 0.0927f
C4187 xaa5.xa3.xb1_0.G CK 0.129f
C4188 xaa5.xa3.xb2_0.G a_26092_62862# 0.00758f
C4189 xaa5.xb1.MN1.G xaa5.xa3.xb2_0.D 0.00217f
C4190 xaa4.xa2.M0.G a_29764_62862# 3.48e-19
C4191 AVDD xaa1.xa3.D 3.18f
C4192 xaa6.xc.XA1.MN0.G xaa6.xd.XA1.MN0.G 0.0191f
C4193 a_29764_58030# a_29764_57678# 0.0109f
C4194 a_36172_58030# xaa6.xf.XA1.MN0.G 0.0408f
C4195 PWRUP_1V8 a_32284_56974# 0.0658f
C4196 AVDD a_34804_56974# 0.00151f
C4197 m2_4468_91484# m3_37748_91804# 0.0138f
C4198 AVDD a_29764_53102# 0.00163f
C4199 xaa6.xd.XA1.MN0.G a_29764_54510# 0.00232f
C4200 xaa6.xc.XA6.MP0.D a_27244_55918# 0.00176f
C4201 xaa6.xg.XA7.MN1.D xaa6.xg.XA3.MN0.D 0.0425f
C4202 xaa6.xg.XA6.MP0.D a_37324_56270# 0.0467f
C4203 xaa6.xf.XA1.MN0.G xaa6.xg.XA3.MP0.D 2.36e-19
C4204 a_34804_56622# xaa6.xf.XA5.MN0.G 6.14e-19
C4205 xaa6.xg.XA3.MP0.D a_37324_54510# 0.0467f
C4206 xaa1.xa4.M0.D m3_4628_102204# 0.0276f
C4207 xaa4.xa2.M0.G m3_13116_54132# 0.0634f
C4208 a_29764_64622# a_29764_64270# 0.0109f
C4209 xaa5.xb3.MP1.D a_28612_64270# 0.0955f
C4210 li_4468_76124# m1_4468_76124# 23f
C4211 xaa1.xa1.M4.D a_n908_59750# 1.21e-19
C4212 xaa3.xa4.MN0.D a_5844_60078# 0.00224f
C4213 a_4692_60430# a_4692_60078# 0.0109f
C4214 PWRUP_1V8 a_32284_58030# 8.58e-19
C4215 AVDD a_34804_58030# 0.00504f
C4216 m2_4468_104924# m3_37668_105244# 0.0138f
C4217 xaa6.xg.XA7.MP1.G a_36172_56270# 0.0985f
C4218 xaa6.xg.XA7.MN1.G a_37324_56270# 0.082f
C4219 xaa6.xf.XA7.MN1.D xaa6.xf.XA5.MN0.G 0.29f
C4220 xaa6.xd.XA7.MP1.G a_28612_55918# 0.0292f
C4221 xaa6.xd.XA7.MN1.G a_27244_55918# 7.1e-20
C4222 a_28612_56622# a_29764_56622# 0.00133f
C4223 xaa6.xc.XA1.MN0.G a_27244_55566# 0.0022f
C4224 xaa1.xa4.M0.D li_4468_116284# 23f
C4225 AVDD xaa6.xg.XA3.MN0.D 0.00913f
C4226 xaa6.xd.XA4.MP0.D a_28612_54862# 0.00176f
C4227 a_27244_55214# a_28612_55214# 8.89e-19
C4228 a_2948_74698# m2_4468_75164# 0.00238f
C4229 xaa1.xa4.M0.D m2_4468_73244# 71.5f
C4230 a_36172_53102# a_37324_53102# 0.00133f
C4231 a_28612_53102# a_28612_52750# 0.0109f
C4232 li_4468_76924# li_4468_76124# 39.3f
C4233 xaa5.xa3.xb2_0.D a_26092_61102# 6.02e-20
C4234 IBPSR_1U a_4692_58142# 1.59e-20
C4235 xaa3.xa1b.MN0.D xaa3.xa2.MN0.D 0.0558f
C4236 xaa4.xa2.M0.G a_11712_59086# 0.0155f
C4237 xaa3.xa5a.MN0.D a_5844_60430# 0.00414f
C4238 AVDD a_29764_62158# 0.00139f
C4239 xaa6.xc.XA7.MN1.G xaa6.xc.XA7.MN2.D 0.0148f
C4240 xaa6.xf.XA1.MN0.G a_34804_56974# 0.00134f
C4241 xaa6.xf.XA7.MN1.D a_36172_56974# 1.31e-19
C4242 xaa6.xd.XA7.MN1.D a_28612_56622# 0.0232f
C4243 xaa6.xc.XA1.MN0.G a_29764_56622# 1.73e-19
C4244 AVDD xaa6.xd.XA5.MN0.G 0.88f
C4245 m2_4468_78044# m3_37748_78364# 0.0138f
C4246 xaa0.xa5.MN2.G a_10092_52750# 3.98e-19
C4247 xaa6.xe.XA5.MN0.G a_32284_55566# 0.0889f
C4248 xaa6.xc.XA7.MP1.G a_27244_53454# 1.07e-19
C4249 xaa6.xc.XA7.MN1.G a_28612_53454# 7.1e-20
C4250 xaa6.xe.XA1.MN0.G a_32284_53102# 0.0711f
C4251 xaa6.xg.XA7.MN1.G a_37324_53806# 0.00785f
C4252 xaa6.xg.XA7.MP1.G a_36172_53806# 0.00375f
C4253 xaa6.xe.XA6.MN0.G xaa6.xe.XA4.MP0.D 0.0357f
C4254 xaa1.xa4.M0.D m1_4468_87644# 67.7f
C4255 xaa4.xa1.M3.D xaa4.xa1.M2.D 0.0488f
C4256 xaa1.xa4.M0.D m3_37668_85084# 0.074f
C4257 xaa1.xa2.M5.D xaa1.xa2.M4.D 0.0488f
C4258 a_4692_62718# a_5844_62718# 0.00133f
C4259 xaa3.xa6.MN0.D xaa3.xa5a.MN0.D 0.187f
C4260 xaa4.xa2.M0.G a_28612_62862# 0.0362f
C4261 xaa5.xb1.MN1.G CK 0.0104f
C4262 xaa5.xa3.xb2_0.G xaa5.xb2_3.MN0.D 0.00946f
C4263 m1_4468_103004# m2_4468_103004# 12.9f
C4264 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN1.D 0.274f
C4265 a_34804_58030# xaa6.xf.XA1.MN0.G 0.00237f
C4266 PWRUP_1V8 a_31132_56974# 0.0768f
C4267 AVDD a_33652_56974# 0.405f
C4268 m2_4468_91484# m3_37668_91804# 0.0138f
C4269 xaa6.xd.XA1.MN0.G a_28612_54510# 1.17e-19
C4270 xaa6.xd.XA7.MN1.D a_29764_54510# 0.072f
C4271 xaa1.xa4.M0.D li_4468_82684# 23f
C4272 PWRUP_1V8 a_26092_53102# 4.2e-19
C4273 xaa6.xg.XA7.MN1.D xaa6.xg.XA3.MN1.G 0.158f
C4274 a_29764_56270# a_31132_56270# 8.89e-19
C4275 xaa6.xe.XA6.MP0.D xaa6.xe.XA6.MN0.G 0.0116f
C4276 xaa6.xg.XA6.MN0.D a_37324_56270# 2.16e-19
C4277 xaa6.xg.XA6.MP0.D a_36172_56270# 2.16e-19
C4278 xaa6.xf.XA1.MN0.G xaa6.xg.XA3.MN0.D 0.00287f
C4279 xaa6.xd.XA7.MN1.G a_29764_54862# 0.0708f
C4280 AVDD a_28612_53102# 0.488f
C4281 xaa6.xd.XA3.MP0.D a_28612_54158# 0.00176f
C4282 a_29764_54510# a_31132_54510# 8.89e-19
C4283 xaa6.xg.XA3.MN0.D a_37324_54510# 2.16e-19
C4284 xaa6.xg.XA3.MP0.D a_36172_54510# 2.16e-19
C4285 xaa1.xa4.M0.D m3_37748_102364# 0.111f
C4286 xaa4.xa2.M0.G m3_13044_54132# 0.106f
C4287 li_4468_110684# li_4468_110524# 7.91f
C4288 xaa3.xa4.MN0.D a_4692_60078# 0.00346f
C4289 a_5844_60430# xaa3.xa3a.MN0.D 0.0658f
C4290 xaa1.xa1.M1.D xaa1.xa1.M0.D 0.0488f
C4291 PWRUP_1V8 a_31132_58030# 0.00223f
C4292 AVDD a_33652_58030# 0.338f
C4293 xaa6.xc.XA7.MN1.D a_27244_55566# 0.00147f
C4294 a_34804_56974# a_34804_56622# 0.0109f
C4295 xaa6.xe.XA7.MN0.D xaa6.xe.XA6.MN0.G 3.13e-19
C4296 xaa6.xc.XA1.MN0.G a_26092_55566# 1.25e-19
C4297 xaa6.xe.XA1.MN0.G xaa6.xf.XA5.MN0.G 0.00881f
C4298 xaa6.xg.XA7.MN1.G a_36172_56270# 0.00344f
C4299 AVDD xaa6.xg.XA3.MN1.G 1.14f
C4300 xaa6.xf.XA5.MN0.G a_34804_54510# 0.00236f
C4301 xaa6.xf.XA4.MN0.D a_34804_55214# 0.0472f
C4302 a_2948_74698# m2_4468_76124# 0.00238f
C4303 xaa1.xa4.M0.D m2_4468_74204# 71.5f
C4304 li_4468_99164# m1_4468_99164# 23f
C4305 a_26092_61806# a_27244_61806# 0.00133f
C4306 xaa5.xb2_0.MN0.D a_29764_61806# 0.126f
C4307 IBPSR_1U xaa3.xa2.MN0.D 3.88e-20
C4308 xaa3.xa5a.MN0.D a_4692_60430# 0.00348f
C4309 xaa5.xa3.xb1_0.D a_28612_61454# 4.81e-19
C4310 AVDD a_28612_62158# 0.352f
C4311 m1_4468_70364# m2_4468_70364# 12.9f
C4312 a_27244_57326# a_28612_57326# 8.89e-19
C4313 xaa6.xf.XA7.MN0.D a_34804_57326# 0.055f
C4314 xaa6.xf.XA7.MN1.D a_34804_56974# 0.0092f
C4315 xaa6.xc.XA1.MN0.G a_28612_56622# 0.00369f
C4316 AVDD xaa6.xc.XA5.MN0.G 0.88f
C4317 m2_4468_78044# m3_37668_78364# 0.0138f
C4318 xaa6.xe.XA7.MN1.D a_32284_53102# 5.24e-20
C4319 xaa6.xe.XA1.MN0.G a_31132_53102# 0.0727f
C4320 xaa6.xe.XA5.MN0.G a_31132_55566# 0.112f
C4321 xaa6.xc.XA7.MP1.G a_26092_53454# 2.78e-19
C4322 xaa6.xc.XA7.MN1.G a_27244_53454# 0.101f
C4323 xaa6.xg.XA7.MN1.G a_36172_53806# 2.31e-19
C4324 xaa6.xe.XA6.MN0.G xaa6.xe.XA4.MN0.D 0.0093f
C4325 xaa6.xe.XA7.MN1.G xaa6.xe.XA1.MN0.D 0.123f
C4326 xaa1.xa4.M0.D m1_4468_88604# 67.7f
C4327 a_29764_53806# a_31132_53806# 8.89e-19
C4328 a_4308_53678# xbb1.xa3.M6.D 5.84e-19
C4329 xaa1.xa4.M0.D m3_4788_85884# 0.0138f
C4330 li_4468_94204# li_4468_93404# 39.3f
C4331 xaa1.xa3.D a_640_61510# 0.0336f
C4332 a_28612_63566# a_28612_63214# 0.0109f
C4333 xaa5.xa3.xb2_0.G a_29764_63214# 0.00375f
C4334 xaa5.xb1.MN1.G a_29764_62862# 0.00532f
C4335 xaa4.xa2.M0.G a_27244_62862# 6.38e-19
C4336 xaa6.xc.XA7.MN1.D xaa6.xd.XA7.MN1.D 0.00435f
C4337 a_28612_58030# a_28612_57678# 0.0109f
C4338 xaa0.xa2a.MN0.D a_244_56270# 6.38e-19
C4339 a_34804_58030# xaa6.xf.XA7.MN1.D 0.0693f
C4340 PWRUP_1V8 a_29764_56974# 0.0755f
C4341 AVDD a_32284_56974# 0.405f
C4342 xaa6.xc.XA1.MN0.G a_29764_54510# 1.02e-19
C4343 xaa6.xd.XA7.MN1.D a_28612_54510# 0.0851f
C4344 xaa6.xf.XA7.MN1.G a_34804_55214# 0.00134f
C4345 xaa6.xg.XA6.MN0.D a_36172_56270# 0.0474f
C4346 xaa6.xe.XA6.MN0.D xaa6.xe.XA6.MN0.G 0.0093f
C4347 xaa6.xf.XA1.MN0.G xaa6.xg.XA3.MN1.G 0.0135f
C4348 xaa6.xd.XA7.MP1.G a_29764_54862# 0.029f
C4349 xaa6.xd.XA7.MN1.G a_28612_54862# 0.00608f
C4350 xaa6.xc.XA6.MN0.D a_26092_55918# 0.00176f
C4351 AVDD a_27244_53102# 0.486f
C4352 xaa6.xg.XA3.MN0.D a_36172_54510# 0.0474f
C4353 xaa6.xg.XA3.MN1.G a_37324_54510# 1.88e-19
C4354 xaa1.xa4.M0.D m3_37668_102364# 0.074f
C4355 xaa4.xa2.M0.G m3_22620_55012# 0.0273f
C4356 a_28612_64622# a_28612_64270# 0.0109f
C4357 xaa1.xa3.D xaa1.xa4.M0.G 0.0605f
C4358 a_4692_60430# xaa3.xa3a.MN0.D 0.0728f
C4359 PWRUP_1V8 a_29764_58030# 0.00667f
C4360 AVDD a_32284_58030# 0.343f
C4361 xaa6.xe.XA7.MP1.G xaa6.xe.XA6.MN0.G 0.524f
C4362 xaa6.xe.XA7.MN1.G xaa6.xf.XA6.MN0.G 3.47e-19
C4363 xaa6.xc.XA7.MN1.D a_26092_55566# 0.00699f
C4364 CK a_36172_54158# 5.04e-20
C4365 a_27244_56622# a_28612_56622# 8.89e-19
C4366 xaa6.xe.XA1.MN0.G xaa6.xe.XA5.MN0.G 0.01f
C4367 xaa1.xa4.M0.D li_4468_117244# 23f
C4368 AVDD xaa6.xf.XA3.MN0.D 0.00913f
C4369 xaa6.xf.XA5.MN0.G a_33652_54510# 0.00224f
C4370 xaa6.xc.XA4.MP0.D a_27244_54862# 0.00176f
C4371 a_26092_55214# a_27244_55214# 0.00133f
C4372 a_2948_74698# m2_4468_77084# 8.4e-19
C4373 xaa1.xa4.M0.D m2_4468_75164# 71.5f
C4374 a_34804_53102# a_36172_53102# 8.89e-19
C4375 a_27244_53102# a_27244_52750# 0.0109f
C4376 li_4468_77084# li_4468_76924# 7.91f
C4377 xaa1.xa2.M2.D PWRUP_1V8 0.00196f
C4378 xaa1.xa2.M1.D a_n908_61510# 5.84e-19
C4379 xaa5.xb2_0.MN0.D a_28612_61806# 0.0878f
C4380 xaa3.xa1b.MN0.D a_4692_58494# 0.00455f
C4381 xaa3.xa5a.MN0.D xaa3.xa4.MN0.D 0.175f
C4382 a_5844_62366# a_5844_60782# 0.00744f
C4383 xaa5.xa3.xb1_0.D a_27244_61454# 0.113f
C4384 AVDD a_27244_62158# 0.384f
C4385 xaa6.xf.XA7.MN1.G a_34804_57326# 0.0797f
C4386 xaa6.xf.XA7.MN0.D a_33652_57326# 0.0525f
C4387 xaa6.xf.XA7.MN1.D a_33652_56974# 0.00166f
C4388 xaa6.xe.XA1.MN0.G a_34804_56974# 0.0677f
C4389 PWRUP_1V8 a_4692_55150# 9.58e-19
C4390 xaa6.xc.XA1.MN0.G a_27244_56622# 0.0022f
C4391 AVDD a_10092_55566# 0.00189f
C4392 xaa6.xe.XA7.MN1.D a_31132_53102# 8.73e-21
C4393 xaa1.xa4.M0.D m1_4468_89564# 67.7f
C4394 xaa6.xc.XA7.MN1.G a_26092_53454# 0.015f
C4395 xaa1.xa4.M0.D m3_4628_85884# 0.0276f
C4396 xaa3.xa6.MN0.D a_5844_62718# 0.0897f
C4397 xaa1.xa3.D a_n908_61510# 3.05e-20
C4398 xaa5.xa3.xb2_0.G a_28612_63214# 0.00581f
C4399 xaa5.xb1.MN1.G a_28612_62862# 9.6e-19
C4400 m1_4468_103964# m2_4468_103964# 12.9f
C4401 xaa0.xa5.MN2.G xaa6.xd.XA7.MN1.D 4.33e-19
C4402 xaa6.xc.XA7.MN1.D xaa6.xc.XA1.MN0.G 0.0209f
C4403 xaa0.xa2a.MN0.D a_n908_56270# 6.26e-20
C4404 a_34804_58030# xaa6.xe.XA1.MN0.G 0.0354f
C4405 a_33652_58030# xaa6.xf.XA7.MN1.D 0.0674f
C4406 PWRUP_1V8 a_28612_56974# 0.0674f
C4407 xaa4.xa2.M0.G a_11712_55918# 0.014f
C4408 AVDD a_31132_56974# 0.00151f
C4409 xaa6.xc.XA1.MN0.G a_28612_54510# 0.00196f
C4410 xaa1.xa4.M0.D li_4468_83644# 23f
C4411 PWRUP_1V8 xaa4.xa1.M0.D 0.00131f
C4412 xaa6.xf.XA7.MP1.G a_34804_55214# 0.096f
C4413 xaa6.xf.XA7.MN1.G a_33652_55214# 0.0745f
C4414 a_28612_56270# a_29764_56270# 0.00133f
C4415 xaa6.xf.XA1.MN0.G xaa6.xf.XA3.MN0.D 0.00303f
C4416 xaa6.xd.XA7.MP1.G a_28612_54862# 0.0986f
C4417 xaa6.xd.XA7.MN1.G a_27244_54862# 7.1e-20
C4418 AVDD a_26092_53102# 0.00171f
C4419 xaa6.xc.XA3.MP0.D a_27244_54158# 0.00176f
C4420 a_28612_54510# a_29764_54510# 0.00133f
C4421 xaa6.xg.XA3.MN1.G a_36172_54510# 0.082f
C4422 xaa1.xa4.M0.D m3_4788_103164# 0.0138f
C4423 xaa4.xa2.M0.G m3_22548_55012# 0.0137f
C4424 li_4468_111484# li_4468_110684# 39.3f
C4425 a_28612_64622# xaa5.xb3.MP1.D 0.0971f
C4426 li_4468_77084# m1_4468_77084# 23f
C4427 xaa3.xa4.MN0.D xaa3.xa3a.MN0.D 0.187f
C4428 PWRUP_1V8 a_28612_58030# 4.25e-19
C4429 AVDD a_31132_58030# 0.00519f
C4430 xaa6.xe.XA7.MN1.G xaa6.xe.XA6.MN0.G 0.329f
C4431 a_33652_56974# a_33652_56622# 0.0109f
C4432 xaa6.xe.XA7.MN1.D xaa6.xe.XA5.MN0.G 0.29f
C4433 xaa3.xa1b.MN0.D xbb1.xa3.M5.D 1.38e-19
C4434 xaa6.xc.XA7.MN1.G a_28612_55918# 7.1e-20
C4435 xaa6.xc.XA7.MP1.G a_27244_55918# 0.0292f
C4436 AVDD xaa6.xf.XA3.MP0.D 0.133f
C4437 xaa6.xf.XA4.MP0.D a_33652_55214# 0.0467f
C4438 xaa1.xa4.M0.D m2_4468_76124# 71.5f
C4439 xaa4.xa2.M0.G xaa4.xa4.M0.D 2.79f
C4440 IBPSR_1U a_4692_58494# 1.59e-20
C4441 xaa5.xa3.xb1_0.D a_26092_61454# 0.0392f
C4442 xaa5.xb2_1.MN0.D PWRUP_1V8 3.2e-20
C4443 AVDD a_26092_62158# 0.00172f
C4444 xaa6.xf.XA7.MN1.G a_33652_57326# 0.00174f
C4445 xaa6.xf.XA7.MP1.G a_34804_57326# 9.02e-20
C4446 xaa6.xc.XA7.MN1.D a_27244_56622# 0.0232f
C4447 xaa6.xe.XA1.MN0.G a_33652_56974# 0.0736f
C4448 PWRUP_1V8 a_5844_55502# 0.0674f
C4449 xaa6.xc.XA1.MN0.G a_26092_56622# 1.25e-19
C4450 a_26092_57326# a_27244_57326# 0.00133f
C4451 AVDD a_5844_55150# 0.443f
C4452 xaa6.xd.XA5.MN0.G a_29764_55566# 0.113f
C4453 xaa6.xd.XA6.MN0.G xaa6.xd.XA4.MN0.D 0.0093f
C4454 xaa1.xa4.M0.D m1_4468_90524# 67.7f
C4455 a_28612_53806# a_29764_53806# 0.00133f
C4456 xaa1.xa4.M0.D m3_37748_86044# 0.111f
C4457 li_4468_94364# li_4468_94204# 7.91f
C4458 xaa3.xa6.MN0.D a_4692_62718# 0.117f
C4459 xaa5.xa3.xb2_0.G a_27244_63214# 0.00829f
C4460 xaa4.xa2.M0.G xaa5.xb2_3.MN0.D 0.174f
C4461 xaa5.xa3.xb1_0.G a_26092_62862# 0.00255f
C4462 xaa0.xa5.MN2.G xaa6.xc.XA1.MN0.G 0.0426f
C4463 a_27244_58030# a_27244_57678# 0.0109f
C4464 xaa0.xa2a.MN0.D xaa0.xa5.MN2.D 7.55e-20
C4465 a_33652_58030# xaa6.xe.XA1.MN0.G 0.0493f
C4466 PWRUP_1V8 a_27244_56974# 0.0658f
C4467 AVDD a_29764_56974# 0.00151f
C4468 xaa6.xc.XA1.MN0.G a_27244_54510# 0.00267f
C4469 PWRUP_1V8 a_37324_53454# 0.0674f
C4470 xaa6.xf.XA7.MP1.G a_33652_55214# 0.027f
C4471 xaa6.xf.XA7.MN1.G a_32284_55214# 7.1e-20
C4472 a_31132_56622# xaa6.xe.XA5.MN0.G 6.14e-19
C4473 xaa6.xf.XA6.MN0.D a_34804_56270# 0.0474f
C4474 xaa6.xd.XA6.MN0.D xaa6.xd.XA6.MN0.G 0.0093f
C4475 xaa6.xf.XA7.MN1.D xaa6.xf.XA3.MN0.D 0.0425f
C4476 xaa6.xf.XA1.MN0.G xaa6.xf.XA3.MP0.D 3.58e-19
C4477 xaa1.xa4.M0.D m3_4628_103164# 0.0276f
C4478 xaa4.xa2.M0.G m3_13116_55188# 0.0634f
C4479 a_28612_64622# a_29764_64622# 0.00133f
C4480 PWRUP_1V8 a_27244_58030# 8.58e-19
C4481 CK a_37324_57678# 5.74e-19
C4482 AVDD a_29764_58030# 0.00504f
C4483 m2_4468_105884# m3_37748_106204# 0.0138f
C4484 a_26092_56622# a_27244_56622# 0.00133f
C4485 xaa6.xf.XA7.MN1.G a_34804_56270# 0.00344f
C4486 xaa1.xa4.M0.D li_4468_118204# 23f
C4487 IBPSR_1U xbb1.xa3.M5.D 0.0485f
C4488 xaa6.xd.XA1.MN0.G xaa6.xe.XA5.MN0.G 0.00856f
C4489 xaa6.xc.XA7.MN1.G a_27244_55918# 0.00733f
C4490 xaa6.xc.XA7.MP1.G a_26092_55918# 0.0294f
C4491 AVDD xaa6.xe.XA3.MP0.D 0.133f
C4492 xaa1.xa4.M0.D m2_4468_77084# 71.5f
C4493 xaa6.xc.XA4.MN0.D a_26092_54862# 0.00176f
C4494 xaa4.xa2.M0.D xaa4.xa1.M5.D 0.00336f
C4495 xaa6.xe.XA5.MN0.G a_32284_54510# 0.00224f
C4496 xbb1.xa3.M5.D a_4308_51918# 8.62e-20
C4497 a_33652_53102# a_34804_53102# 0.00133f
C4498 a_26092_53102# a_26092_52750# 0.0109f
C4499 li_4468_100124# m1_4468_100124# 23f
C4500 li_4468_77884# li_4468_77084# 39.3f
C4501 a_4692_62366# a_4692_60782# 0.00744f
C4502 xaa4.xa2.M0.G a_11712_60670# 0.0119f
C4503 a_29764_62158# a_29764_61806# 0.0109f
C4504 xaa5.xa3.xc2a.D a_27244_61806# 0.0467f
C4505 xaa5.xa3.xb2_0.D xaa5.xa3.xc1a.D 0.0801f
C4506 xaa1.xa2.M2.D xaa1.xa1.M8.D 0.00181f
C4507 m1_4468_71324# m2_4468_71324# 12.9f
C4508 xaa6.xf.XA7.MP1.G a_33652_57326# 0.0948f
C4509 PWRUP_1V8 a_4692_55502# 0.069f
C4510 xaa6.xc.XA7.MN1.D a_26092_56622# 0.0377f
C4511 xaa0.xa5.MN2.G a_27244_56622# 0.00119f
C4512 xaa6.xe.XA1.MN0.G a_32284_56974# 0.00218f
C4513 AVDD a_4692_55150# 0.00527f
C4514 xaa6.xd.XA7.MN1.G xaa6.xd.XA1.MN0.D 0.123f
C4515 xaa6.xd.XA5.MN0.G a_28612_55566# 0.0873f
C4516 xaa6.xd.XA6.MN0.G xaa6.xd.XA4.MP0.D 0.0357f
C4517 xaa6.xd.XA1.MN0.G a_29764_53102# 0.0721f
C4518 xaa1.xa4.M0.D m1_4468_91484# 67.7f
C4519 xaa6.xf.XA7.MN1.G a_34804_53806# 0.115f
C4520 xaa1.xa4.M0.D m3_37668_86044# 0.074f
C4521 a_5844_63070# a_5844_62718# 0.0109f
C4522 xaa5.xa3.xb2_0.G a_26092_63214# 0.0112f
C4523 xaa4.xa2.M0.G a_29764_63214# 3.48e-19
C4524 m1_4468_104924# m2_4468_104924# 12.9f
C4525 a_11712_59086# a_11712_57502# 0.00223f
C4526 xaa0.xa2a.MN0.D xaa0.xa5.MN0.D 0.0021f
C4527 xaa0.xa5.MN2.G xaa6.xc.XA7.MN1.D 0.248f
C4528 a_32284_58030# xaa6.xe.XA1.MN0.G 0.0026f
C4529 PWRUP_1V8 a_26092_56974# 0.077f
C4530 AVDD a_28612_56974# 0.405f
C4531 m2_4468_92444# m3_37748_92764# 0.0138f
C4532 xaa1.xa4.M0.D li_4468_84604# 23f
C4533 xaa6.xc.XA1.MN0.G a_26092_54510# 6.72e-19
C4534 PWRUP_1V8 a_36172_53454# 0.0689f
C4535 a_27244_56270# a_28612_56270# 8.89e-19
C4536 xaa6.xd.XA6.MP0.D xaa6.xd.XA6.MN0.G 0.0116f
C4537 xaa6.xf.XA6.MP0.D a_34804_56270# 2.16e-19
C4538 xaa6.xf.XA6.MN0.D a_33652_56270# 2.16e-19
C4539 xaa6.xc.XA7.MN1.D a_27244_54510# 0.0836f
C4540 xaa6.xf.XA7.MN1.D xaa6.xf.XA3.MP0.D 0.0844f
C4541 xaa6.xe.XA1.MN0.G xaa6.xf.XA3.MN0.D 3.2e-19
C4542 AVDD xaa4.xa1.M0.D 0.00461f
C4543 m3_22620_52900# AVSS 0.174f
C4544 m3_22548_52900# AVSS 0.0651f $ **FLOATING
C4545 m3_13116_53076# AVSS 0.0153f $ **FLOATING
C4546 m3_13044_53076# AVSS 0.0162f
C4547 m3_22620_53956# AVSS 0.174f
C4548 m3_22548_53956# AVSS 0.0651f $ **FLOATING
C4549 m3_13116_54132# AVSS 0.0153f $ **FLOATING
C4550 m3_13044_54132# AVSS 0.0162f
C4551 m3_22620_55012# AVSS 0.174f
C4552 m3_22548_55012# AVSS 0.0651f $ **FLOATING
C4553 m3_13116_55188# AVSS 0.0153f $ **FLOATING
C4554 m3_13044_55188# AVSS 0.0162f
C4555 m3_22620_56068# AVSS 0.174f
C4556 m3_22548_56068# AVSS 0.0651f $ **FLOATING
C4557 m3_13116_56244# AVSS 0.0153f $ **FLOATING
C4558 m3_13044_56244# AVSS 0.0162f
C4559 m3_22620_57124# AVSS 0.174f
C4560 m3_22548_57124# AVSS 0.0651f $ **FLOATING
C4561 m3_13116_57300# AVSS 0.0153f $ **FLOATING
C4562 m3_13044_57300# AVSS 0.0162f
C4563 m3_22620_58180# AVSS 0.174f
C4564 m3_22548_58180# AVSS 0.0651f $ **FLOATING
C4565 m3_13116_58356# AVSS 0.0153f $ **FLOATING
C4566 m3_13044_58356# AVSS 0.0162f
C4567 m3_22620_59236# AVSS 0.174f
C4568 m3_22548_59236# AVSS 0.0651f $ **FLOATING
C4569 m3_13116_59412# AVSS 0.0153f $ **FLOATING
C4570 m3_13044_59412# AVSS 0.0162f
C4571 m3_22620_60292# AVSS 0.174f
C4572 m3_22548_60292# AVSS 0.0651f $ **FLOATING
C4573 m3_13116_60468# AVSS 0.0153f $ **FLOATING
C4574 m3_13044_60468# AVSS 0.0162f
C4575 m3_22620_61348# AVSS 0.174f
C4576 m3_22548_61348# AVSS 0.0651f $ **FLOATING
C4577 m3_13116_61524# AVSS 0.0153f $ **FLOATING
C4578 m3_13044_61524# AVSS 0.0162f
C4579 m3_4788_69564# AVSS 0.0757f $ **FLOATING
C4580 m3_4628_69564# AVSS 0.189f
C4581 m3_37748_69724# AVSS 0.00253f
C4582 m3_37668_69724# AVSS 0.00169f $ **FLOATING
C4583 m3_4788_70524# AVSS 0.0757f $ **FLOATING
C4584 m3_4628_70524# AVSS 0.189f
C4585 m3_37748_70684# AVSS 0.00253f
C4586 m3_37668_70684# AVSS 0.00169f $ **FLOATING
C4587 m3_4788_71484# AVSS 0.0757f $ **FLOATING
C4588 m3_4628_71484# AVSS 0.189f
C4589 m3_37748_71644# AVSS 0.00253f
C4590 m3_37668_71644# AVSS 0.00169f $ **FLOATING
C4591 m3_4788_72444# AVSS 0.0757f $ **FLOATING
C4592 m3_4628_72444# AVSS 0.189f
C4593 m3_37748_72604# AVSS 0.00253f
C4594 m3_37668_72604# AVSS 0.00169f $ **FLOATING
C4595 m3_4788_73404# AVSS 0.0757f $ **FLOATING
C4596 m3_4628_73404# AVSS 0.189f
C4597 m3_37748_73564# AVSS 0.00253f
C4598 m3_37668_73564# AVSS 0.00169f $ **FLOATING
C4599 m3_4788_74364# AVSS 0.0757f $ **FLOATING
C4600 m3_4628_74364# AVSS 0.189f
C4601 m3_37748_74524# AVSS 0.00253f
C4602 m3_37668_74524# AVSS 0.00169f $ **FLOATING
C4603 m3_4788_75324# AVSS 0.0757f $ **FLOATING
C4604 m3_4628_75324# AVSS 0.189f
C4605 m3_37748_75484# AVSS 0.00253f
C4606 m3_37668_75484# AVSS 0.00169f $ **FLOATING
C4607 m3_4788_76284# AVSS 0.0757f $ **FLOATING
C4608 m3_4628_76284# AVSS 0.189f
C4609 m3_37748_76444# AVSS 0.00253f
C4610 m3_37668_76444# AVSS 0.00169f $ **FLOATING
C4611 m3_4788_77244# AVSS 0.0757f $ **FLOATING
C4612 m3_4628_77244# AVSS 0.189f
C4613 m3_37748_77404# AVSS 0.00253f
C4614 m3_37668_77404# AVSS 0.00169f $ **FLOATING
C4615 m3_4788_78204# AVSS 0.0757f $ **FLOATING
C4616 m3_4628_78204# AVSS 0.189f
C4617 m3_37748_78364# AVSS 0.00253f
C4618 m3_37668_78364# AVSS 0.00169f $ **FLOATING
C4619 m3_4788_79164# AVSS 0.0757f $ **FLOATING
C4620 m3_4628_79164# AVSS 0.189f
C4621 m3_37748_79324# AVSS 0.00253f
C4622 m3_37668_79324# AVSS 0.00169f $ **FLOATING
C4623 m3_4788_80124# AVSS 0.0757f $ **FLOATING
C4624 m3_4628_80124# AVSS 0.189f
C4625 m3_37748_80284# AVSS 0.00253f
C4626 m3_37668_80284# AVSS 0.00169f $ **FLOATING
C4627 m3_4788_81084# AVSS 0.0757f $ **FLOATING
C4628 m3_4628_81084# AVSS 0.189f
C4629 m3_37748_81244# AVSS 0.00253f
C4630 m3_37668_81244# AVSS 0.00169f $ **FLOATING
C4631 m3_4788_82044# AVSS 0.0757f $ **FLOATING
C4632 m3_4628_82044# AVSS 0.189f
C4633 m3_37748_82204# AVSS 0.00253f
C4634 m3_37668_82204# AVSS 0.00169f $ **FLOATING
C4635 m3_4788_83004# AVSS 0.0757f $ **FLOATING
C4636 m3_4628_83004# AVSS 0.189f
C4637 m3_37748_83164# AVSS 0.00253f
C4638 m3_37668_83164# AVSS 0.00169f $ **FLOATING
C4639 m3_4788_83964# AVSS 0.0757f $ **FLOATING
C4640 m3_4628_83964# AVSS 0.189f
C4641 m3_37748_84124# AVSS 0.00253f
C4642 m3_37668_84124# AVSS 0.00169f $ **FLOATING
C4643 m3_4788_84924# AVSS 0.0757f $ **FLOATING
C4644 m3_4628_84924# AVSS 0.189f
C4645 m3_37748_85084# AVSS 0.00253f
C4646 m3_37668_85084# AVSS 0.00169f $ **FLOATING
C4647 m3_4788_85884# AVSS 0.0757f $ **FLOATING
C4648 m3_4628_85884# AVSS 0.189f
C4649 m3_37748_86044# AVSS 0.00253f
C4650 m3_37668_86044# AVSS 0.00169f $ **FLOATING
C4651 m3_4788_86844# AVSS 0.0757f $ **FLOATING
C4652 m3_4628_86844# AVSS 0.189f
C4653 m3_37748_87004# AVSS 0.00253f
C4654 m3_37668_87004# AVSS 0.00169f $ **FLOATING
C4655 m3_4788_87804# AVSS 0.0757f $ **FLOATING
C4656 m3_4628_87804# AVSS 0.189f
C4657 m3_37748_87964# AVSS 0.00253f
C4658 m3_37668_87964# AVSS 0.00169f $ **FLOATING
C4659 m3_4788_88764# AVSS 0.0757f $ **FLOATING
C4660 m3_4628_88764# AVSS 0.189f
C4661 m3_37748_88924# AVSS 0.00253f
C4662 m3_37668_88924# AVSS 0.00169f $ **FLOATING
C4663 m3_4788_89724# AVSS 0.0757f $ **FLOATING
C4664 m3_4628_89724# AVSS 0.189f
C4665 m3_37748_89884# AVSS 0.00253f
C4666 m3_37668_89884# AVSS 0.00169f $ **FLOATING
C4667 m3_4788_90684# AVSS 0.0757f $ **FLOATING
C4668 m3_4628_90684# AVSS 0.189f
C4669 m3_37748_90844# AVSS 0.00253f
C4670 m3_37668_90844# AVSS 0.00169f $ **FLOATING
C4671 m3_4788_91644# AVSS 0.0757f $ **FLOATING
C4672 m3_4628_91644# AVSS 0.189f
C4673 m3_37748_91804# AVSS 0.00253f
C4674 m3_37668_91804# AVSS 0.00169f $ **FLOATING
C4675 m3_4788_92604# AVSS 0.0757f $ **FLOATING
C4676 m3_4628_92604# AVSS 0.189f
C4677 m3_37748_92764# AVSS 0.00253f
C4678 m3_37668_92764# AVSS 0.00169f $ **FLOATING
C4679 m3_4788_93564# AVSS 0.0757f $ **FLOATING
C4680 m3_4628_93564# AVSS 0.189f
C4681 m3_37748_93724# AVSS 0.00253f
C4682 m3_37668_93724# AVSS 0.00169f $ **FLOATING
C4683 m3_4788_94524# AVSS 0.0757f $ **FLOATING
C4684 m3_4628_94524# AVSS 0.189f
C4685 m3_37748_94684# AVSS 0.00253f
C4686 m3_37668_94684# AVSS 0.00169f $ **FLOATING
C4687 m3_4788_95484# AVSS 0.0757f $ **FLOATING
C4688 m3_4628_95484# AVSS 0.189f
C4689 m3_37748_95644# AVSS 0.00253f
C4690 m3_37668_95644# AVSS 0.00169f $ **FLOATING
C4691 m3_4788_96444# AVSS 0.0757f $ **FLOATING
C4692 m3_4628_96444# AVSS 0.189f
C4693 m3_37748_96604# AVSS 0.00253f
C4694 m3_37668_96604# AVSS 0.00169f $ **FLOATING
C4695 m3_4788_97404# AVSS 0.0757f $ **FLOATING
C4696 m3_4628_97404# AVSS 0.189f
C4697 m3_37748_97564# AVSS 0.00253f
C4698 m3_37668_97564# AVSS 0.00169f $ **FLOATING
C4699 m3_4788_98364# AVSS 0.0757f $ **FLOATING
C4700 m3_4628_98364# AVSS 0.189f
C4701 m3_37748_98524# AVSS 0.00253f
C4702 m3_37668_98524# AVSS 0.00169f $ **FLOATING
C4703 m3_4788_99324# AVSS 0.0757f $ **FLOATING
C4704 m3_4628_99324# AVSS 0.189f
C4705 m3_37748_99484# AVSS 0.00253f
C4706 m3_37668_99484# AVSS 0.00169f $ **FLOATING
C4707 m3_4788_100284# AVSS 0.0757f $ **FLOATING
C4708 m3_4628_100284# AVSS 0.189f
C4709 m3_37748_100444# AVSS 0.00253f
C4710 m3_37668_100444# AVSS 0.00169f $ **FLOATING
C4711 m3_4788_101244# AVSS 0.0757f $ **FLOATING
C4712 m3_4628_101244# AVSS 0.189f
C4713 m3_37748_101404# AVSS 0.00253f
C4714 m3_37668_101404# AVSS 0.00169f $ **FLOATING
C4715 m3_4788_102204# AVSS 0.0757f $ **FLOATING
C4716 m3_4628_102204# AVSS 0.189f
C4717 m3_37748_102364# AVSS 0.00253f
C4718 m3_37668_102364# AVSS 0.00169f $ **FLOATING
C4719 m3_4788_103164# AVSS 0.0757f $ **FLOATING
C4720 m3_4628_103164# AVSS 0.189f
C4721 m3_37748_103324# AVSS 0.00253f
C4722 m3_37668_103324# AVSS 0.00169f $ **FLOATING
C4723 m3_4788_104124# AVSS 0.0757f $ **FLOATING
C4724 m3_4628_104124# AVSS 0.189f
C4725 m3_37748_104284# AVSS 0.00253f
C4726 m3_37668_104284# AVSS 0.00169f $ **FLOATING
C4727 m3_4788_105084# AVSS 0.0757f $ **FLOATING
C4728 m3_4628_105084# AVSS 0.189f
C4729 m3_37748_105244# AVSS 0.00253f
C4730 m3_37668_105244# AVSS 0.00169f $ **FLOATING
C4731 m3_4788_106044# AVSS 0.0757f $ **FLOATING
C4732 m3_4628_106044# AVSS 0.189f
C4733 m3_37748_106204# AVSS 0.00253f
C4734 m3_37668_106204# AVSS 0.00169f $ **FLOATING
C4735 m3_4788_107004# AVSS 0.0757f $ **FLOATING
C4736 m3_4628_107004# AVSS 0.189f
C4737 m3_37748_107164# AVSS 0.00253f
C4738 m3_37668_107164# AVSS 0.00169f $ **FLOATING
C4739 m3_4788_107964# AVSS 0.0757f $ **FLOATING
C4740 m3_4628_107964# AVSS 0.189f
C4741 m3_37748_108124# AVSS 0.00253f
C4742 m3_37668_108124# AVSS 0.00169f $ **FLOATING
C4743 m3_4788_108924# AVSS 0.0757f $ **FLOATING
C4744 m3_4628_108924# AVSS 0.189f
C4745 m3_37748_109084# AVSS 0.00253f
C4746 m3_37668_109084# AVSS 0.00169f $ **FLOATING
C4747 m3_4788_109884# AVSS 0.0757f $ **FLOATING
C4748 m3_4628_109884# AVSS 0.189f
C4749 m3_37748_110044# AVSS 0.00253f
C4750 m3_37668_110044# AVSS 0.00169f $ **FLOATING
C4751 m3_4788_110844# AVSS 0.0757f $ **FLOATING
C4752 m3_4628_110844# AVSS 0.189f
C4753 m3_37748_111004# AVSS 0.00253f
C4754 m3_37668_111004# AVSS 0.00169f $ **FLOATING
C4755 m3_4788_111804# AVSS 0.0757f $ **FLOATING
C4756 m3_4628_111804# AVSS 0.189f
C4757 m3_37748_111964# AVSS 0.00253f
C4758 m3_37668_111964# AVSS 0.00169f $ **FLOATING
C4759 m3_4788_112764# AVSS 0.0757f $ **FLOATING
C4760 m3_4628_112764# AVSS 0.189f
C4761 m3_37748_112924# AVSS 0.00253f
C4762 m3_37668_112924# AVSS 0.00169f $ **FLOATING
C4763 m3_4788_113724# AVSS 0.0757f $ **FLOATING
C4764 m3_4628_113724# AVSS 0.189f
C4765 m3_37748_113884# AVSS 0.00253f
C4766 m3_37668_113884# AVSS 0.00169f $ **FLOATING
C4767 m3_4788_114684# AVSS 0.0757f $ **FLOATING
C4768 m3_4628_114684# AVSS 0.189f
C4769 m3_37748_114844# AVSS 0.00253f
C4770 m3_37668_114844# AVSS 0.00169f $ **FLOATING
C4771 m3_4788_115644# AVSS 0.0757f $ **FLOATING
C4772 m3_4628_115644# AVSS 0.189f
C4773 m3_37748_115804# AVSS 0.00253f
C4774 m3_37668_115804# AVSS 0.00169f $ **FLOATING
C4775 m3_4788_116604# AVSS 0.0757f $ **FLOATING
C4776 m3_4628_116604# AVSS 0.189f
C4777 m3_37748_116764# AVSS 0.00253f
C4778 m3_37668_116764# AVSS 0.00169f $ **FLOATING
C4779 m3_4788_117564# AVSS 0.0757f $ **FLOATING
C4780 m3_4628_117564# AVSS 0.189f
C4781 m3_37748_117724# AVSS 0.00253f
C4782 m3_37668_117724# AVSS 0.00169f $ **FLOATING
C4783 m2_4468_69404# AVSS 25.9f $ **FLOATING
C4784 m2_4468_70364# AVSS 20f $ **FLOATING
C4785 m2_4468_71324# AVSS 20f $ **FLOATING
C4786 m2_4468_72284# AVSS 20f $ **FLOATING
C4787 m2_4468_73244# AVSS 20f $ **FLOATING
C4788 m2_4468_74204# AVSS 20f $ **FLOATING
C4789 m2_4468_75164# AVSS 20f $ **FLOATING
C4790 m2_4468_76124# AVSS 20f $ **FLOATING
C4791 m2_4468_77084# AVSS 20f $ **FLOATING
C4792 m2_4468_78044# AVSS 20f $ **FLOATING
C4793 m2_4468_79004# AVSS 20f $ **FLOATING
C4794 m2_4468_79964# AVSS 20f $ **FLOATING
C4795 m2_4468_80924# AVSS 20f $ **FLOATING
C4796 m2_4468_81884# AVSS 20f $ **FLOATING
C4797 m2_4468_82844# AVSS 20f $ **FLOATING
C4798 m2_4468_83804# AVSS 20f $ **FLOATING
C4799 m2_4468_84764# AVSS 20f $ **FLOATING
C4800 m2_4468_85724# AVSS 20f $ **FLOATING
C4801 m2_4468_86684# AVSS 20f $ **FLOATING
C4802 m2_4468_87644# AVSS 20f $ **FLOATING
C4803 m2_4468_88604# AVSS 20f $ **FLOATING
C4804 m2_4468_89564# AVSS 20f $ **FLOATING
C4805 m2_4468_90524# AVSS 20f $ **FLOATING
C4806 m2_4468_91484# AVSS 20f $ **FLOATING
C4807 m2_4468_92444# AVSS 20f $ **FLOATING
C4808 m2_4468_93404# AVSS 20f $ **FLOATING
C4809 m2_4468_94364# AVSS 20f $ **FLOATING
C4810 m2_4468_95324# AVSS 20f $ **FLOATING
C4811 m2_4468_96284# AVSS 20f $ **FLOATING
C4812 m2_4468_97244# AVSS 20f $ **FLOATING
C4813 m2_4468_98204# AVSS 20f $ **FLOATING
C4814 m2_4468_99164# AVSS 20f $ **FLOATING
C4815 m2_4468_100124# AVSS 20f $ **FLOATING
C4816 m2_4468_101084# AVSS 20f $ **FLOATING
C4817 m2_4468_102044# AVSS 20f $ **FLOATING
C4818 m2_4468_103004# AVSS 20f $ **FLOATING
C4819 m2_4468_103964# AVSS 20f $ **FLOATING
C4820 m2_4468_104924# AVSS 20f $ **FLOATING
C4821 m2_4468_105884# AVSS 20f $ **FLOATING
C4822 m2_4468_106844# AVSS 20f $ **FLOATING
C4823 m2_4468_107804# AVSS 20f $ **FLOATING
C4824 m2_4468_108764# AVSS 20f $ **FLOATING
C4825 m2_4468_109724# AVSS 20f $ **FLOATING
C4826 m2_4468_110684# AVSS 20f $ **FLOATING
C4827 m2_4468_111644# AVSS 20f $ **FLOATING
C4828 m2_4468_112604# AVSS 20f $ **FLOATING
C4829 m2_4468_113564# AVSS 20f $ **FLOATING
C4830 m2_4468_114524# AVSS 20f $ **FLOATING
C4831 m2_4468_115484# AVSS 20f $ **FLOATING
C4832 m2_4468_116444# AVSS 20f $ **FLOATING
C4833 m2_4468_117404# AVSS 20f $ **FLOATING
C4834 m1_37504_55818# AVSS 0.014f $ **FLOATING
C4835 m1_37504_57930# AVSS 0.0621f $ **FLOATING
C4836 m1_4468_69404# AVSS 12.2f $ **FLOATING
C4837 m1_4468_70204# AVSS 5.5f $ **FLOATING
C4838 m1_4468_70364# AVSS 5.51f $ **FLOATING
C4839 m1_4468_71164# AVSS 5.5f $ **FLOATING
C4840 m1_4468_71324# AVSS 5.51f $ **FLOATING
C4841 m1_4468_72124# AVSS 5.5f $ **FLOATING
C4842 m1_4468_72284# AVSS 5.51f $ **FLOATING
C4843 m1_4468_73244# AVSS 5.51f $ **FLOATING
C4844 m1_4468_74204# AVSS 5.51f $ **FLOATING
C4845 m1_4468_75164# AVSS 5.51f $ **FLOATING
C4846 m1_4468_76124# AVSS 5.51f $ **FLOATING
C4847 m1_4468_77084# AVSS 5.51f $ **FLOATING
C4848 m1_4468_78044# AVSS 5.51f $ **FLOATING
C4849 m1_4468_79004# AVSS 5.51f $ **FLOATING
C4850 m1_4468_79964# AVSS 5.51f $ **FLOATING
C4851 m1_4468_80924# AVSS 5.51f $ **FLOATING
C4852 m1_4468_81884# AVSS 5.51f $ **FLOATING
C4853 m1_4468_82844# AVSS 5.51f $ **FLOATING
C4854 m1_4468_83804# AVSS 5.51f $ **FLOATING
C4855 m1_4468_84764# AVSS 5.51f $ **FLOATING
C4856 m1_4468_85724# AVSS 5.51f $ **FLOATING
C4857 m1_4468_86684# AVSS 5.51f $ **FLOATING
C4858 m1_4468_87644# AVSS 5.51f $ **FLOATING
C4859 m1_4468_88604# AVSS 5.51f $ **FLOATING
C4860 m1_4468_89564# AVSS 5.51f $ **FLOATING
C4861 m1_4468_90524# AVSS 5.51f $ **FLOATING
C4862 m1_4468_91484# AVSS 5.51f $ **FLOATING
C4863 m1_4468_92444# AVSS 5.51f $ **FLOATING
C4864 m1_4468_93404# AVSS 5.51f $ **FLOATING
C4865 m1_4468_94364# AVSS 5.51f $ **FLOATING
C4866 m1_4468_95324# AVSS 5.51f $ **FLOATING
C4867 m1_4468_96284# AVSS 5.51f $ **FLOATING
C4868 m1_4468_97244# AVSS 5.51f $ **FLOATING
C4869 m1_4468_98204# AVSS 5.51f $ **FLOATING
C4870 m1_4468_99164# AVSS 5.51f $ **FLOATING
C4871 m1_4468_100124# AVSS 5.51f $ **FLOATING
C4872 m1_4468_101084# AVSS 5.51f $ **FLOATING
C4873 m1_4468_102044# AVSS 5.51f $ **FLOATING
C4874 m1_4468_103004# AVSS 5.51f $ **FLOATING
C4875 m1_4468_103964# AVSS 5.51f $ **FLOATING
C4876 m1_4468_104924# AVSS 5.51f $ **FLOATING
C4877 m1_4468_105884# AVSS 5.51f $ **FLOATING
C4878 m1_4468_106844# AVSS 5.51f $ **FLOATING
C4879 m1_4468_107804# AVSS 5.51f $ **FLOATING
C4880 m1_4468_108764# AVSS 5.51f $ **FLOATING
C4881 m1_4468_109724# AVSS 5.51f $ **FLOATING
C4882 m1_4468_110684# AVSS 5.51f $ **FLOATING
C4883 m1_4468_111644# AVSS 5.51f $ **FLOATING
C4884 m1_4468_112604# AVSS 5.51f $ **FLOATING
C4885 m1_4468_113564# AVSS 5.51f $ **FLOATING
C4886 m1_4468_114524# AVSS 5.51f $ **FLOATING
C4887 m1_4468_115484# AVSS 5.51f $ **FLOATING
C4888 m1_4468_116444# AVSS 5.51f $ **FLOATING
C4889 m1_4468_117404# AVSS 5.51f $ **FLOATING
C4890 li_4980_56708# AVSS 0.0438f $ **FLOATING
C4891 li_4836_56708# AVSS 0.115f
C4892 li_6204_57236# AVSS 0.0382f
C4893 li_6132_57236# AVSS 0.0117f $ **FLOATING
C4894 li_4980_58996# AVSS 0.0438f $ **FLOATING
C4895 li_4836_58996# AVSS 0.115f
C4896 li_6204_59524# AVSS 0.0382f
C4897 li_6132_59524# AVSS 0.0117f $ **FLOATING
C4898 li_4980_61284# AVSS 0.0438f $ **FLOATING
C4899 li_4836_61284# AVSS 0.115f
C4900 li_6204_61812# AVSS 0.0382f
C4901 li_6132_61812# AVSS 0.0117f $ **FLOATING
C4902 li_4468_69404# AVSS 22f $ **FLOATING
C4903 li_4468_70204# AVSS 15.2f $ **FLOATING
C4904 li_4468_70364# AVSS 15.2f $ **FLOATING
C4905 li_4468_71164# AVSS 15.2f $ **FLOATING
C4906 li_4468_71324# AVSS 15.2f $ **FLOATING
C4907 li_4468_72124# AVSS 15.2f $ **FLOATING
C4908 li_4468_72284# AVSS 15.2f $ **FLOATING
C4909 li_4468_73084# AVSS 15.2f $ **FLOATING
C4910 li_4468_73244# AVSS 15.2f $ **FLOATING
C4911 li_4468_74044# AVSS 15.2f $ **FLOATING
C4912 li_4468_74204# AVSS 15.2f $ **FLOATING
C4913 li_4468_75004# AVSS 15.2f $ **FLOATING
C4914 li_4468_75164# AVSS 15.2f $ **FLOATING
C4915 li_4468_75964# AVSS 15.2f $ **FLOATING
C4916 li_4468_76124# AVSS 15.2f $ **FLOATING
C4917 li_4468_76924# AVSS 15.2f $ **FLOATING
C4918 li_4468_77084# AVSS 15.2f $ **FLOATING
C4919 li_4468_77884# AVSS 15.2f $ **FLOATING
C4920 li_4468_78044# AVSS 15.2f $ **FLOATING
C4921 li_4468_78844# AVSS 15.2f $ **FLOATING
C4922 li_4468_79004# AVSS 15.2f $ **FLOATING
C4923 li_4468_79804# AVSS 15.2f $ **FLOATING
C4924 li_4468_79964# AVSS 15.2f $ **FLOATING
C4925 li_4468_80764# AVSS 15.2f $ **FLOATING
C4926 li_4468_80924# AVSS 15.2f $ **FLOATING
C4927 li_4468_81724# AVSS 15.2f $ **FLOATING
C4928 li_4468_81884# AVSS 15.2f $ **FLOATING
C4929 li_4468_82684# AVSS 15.2f $ **FLOATING
C4930 li_4468_82844# AVSS 15.2f $ **FLOATING
C4931 li_4468_83644# AVSS 15.2f $ **FLOATING
C4932 li_4468_83804# AVSS 15.2f $ **FLOATING
C4933 li_4468_84604# AVSS 15.2f $ **FLOATING
C4934 li_4468_84764# AVSS 15.2f $ **FLOATING
C4935 li_4468_85564# AVSS 15.2f $ **FLOATING
C4936 li_4468_85724# AVSS 15.2f $ **FLOATING
C4937 li_4468_86524# AVSS 15.2f $ **FLOATING
C4938 li_4468_86684# AVSS 15.2f $ **FLOATING
C4939 li_4468_87484# AVSS 15.2f $ **FLOATING
C4940 li_4468_87644# AVSS 15.2f $ **FLOATING
C4941 li_4468_88444# AVSS 15.2f $ **FLOATING
C4942 li_4468_88604# AVSS 15.2f $ **FLOATING
C4943 li_4468_89404# AVSS 15.2f $ **FLOATING
C4944 li_4468_89564# AVSS 15.2f $ **FLOATING
C4945 li_4468_90364# AVSS 15.2f $ **FLOATING
C4946 li_4468_90524# AVSS 15.2f $ **FLOATING
C4947 li_4468_91324# AVSS 15.2f $ **FLOATING
C4948 li_4468_91484# AVSS 15.2f $ **FLOATING
C4949 li_4468_92284# AVSS 15.2f $ **FLOATING
C4950 li_4468_92444# AVSS 15.2f $ **FLOATING
C4951 li_4468_93244# AVSS 15.2f $ **FLOATING
C4952 li_4468_93404# AVSS 15.2f $ **FLOATING
C4953 li_4468_94204# AVSS 15.2f $ **FLOATING
C4954 li_4468_94364# AVSS 15.2f $ **FLOATING
C4955 li_4468_95164# AVSS 15.2f $ **FLOATING
C4956 li_4468_95324# AVSS 15.2f $ **FLOATING
C4957 li_4468_96124# AVSS 15.2f $ **FLOATING
C4958 li_4468_96284# AVSS 15.2f $ **FLOATING
C4959 li_4468_97084# AVSS 15.2f $ **FLOATING
C4960 li_4468_97244# AVSS 15.2f $ **FLOATING
C4961 li_4468_98044# AVSS 15.2f $ **FLOATING
C4962 li_4468_98204# AVSS 15.2f $ **FLOATING
C4963 li_4468_99004# AVSS 15.2f $ **FLOATING
C4964 li_4468_99164# AVSS 15.2f $ **FLOATING
C4965 li_4468_99964# AVSS 15.2f $ **FLOATING
C4966 li_4468_100124# AVSS 15.2f $ **FLOATING
C4967 li_4468_100924# AVSS 15.2f $ **FLOATING
C4968 li_4468_101084# AVSS 15.2f $ **FLOATING
C4969 li_4468_101884# AVSS 15.2f $ **FLOATING
C4970 li_4468_102044# AVSS 15.2f $ **FLOATING
C4971 li_4468_102844# AVSS 15.2f $ **FLOATING
C4972 li_4468_103004# AVSS 15.2f $ **FLOATING
C4973 li_4468_103804# AVSS 15.2f $ **FLOATING
C4974 li_4468_103964# AVSS 15.2f $ **FLOATING
C4975 li_4468_104764# AVSS 15.2f $ **FLOATING
C4976 li_4468_104924# AVSS 15.2f $ **FLOATING
C4977 li_4468_105724# AVSS 15.2f $ **FLOATING
C4978 li_4468_105884# AVSS 15.2f $ **FLOATING
C4979 li_4468_106684# AVSS 15.2f $ **FLOATING
C4980 li_4468_106844# AVSS 15.2f $ **FLOATING
C4981 li_4468_107644# AVSS 15.2f $ **FLOATING
C4982 li_4468_107804# AVSS 15.2f $ **FLOATING
C4983 li_4468_108604# AVSS 15.2f $ **FLOATING
C4984 li_4468_108764# AVSS 15.2f $ **FLOATING
C4985 li_4468_109564# AVSS 15.2f $ **FLOATING
C4986 li_4468_109724# AVSS 15.2f $ **FLOATING
C4987 li_4468_110524# AVSS 15.2f $ **FLOATING
C4988 li_4468_110684# AVSS 15.2f $ **FLOATING
C4989 li_4468_111484# AVSS 15.2f $ **FLOATING
C4990 li_4468_111644# AVSS 15.2f $ **FLOATING
C4991 li_4468_112444# AVSS 15.2f $ **FLOATING
C4992 li_4468_112604# AVSS 15.2f $ **FLOATING
C4993 li_4468_113404# AVSS 15.2f $ **FLOATING
C4994 li_4468_113564# AVSS 15.2f $ **FLOATING
C4995 li_4468_114364# AVSS 15.2f $ **FLOATING
C4996 li_4468_114524# AVSS 15.2f $ **FLOATING
C4997 li_4468_115324# AVSS 15.2f $ **FLOATING
C4998 li_4468_115484# AVSS 15.2f $ **FLOATING
C4999 li_4468_116284# AVSS 15.2f $ **FLOATING
C5000 li_4468_116444# AVSS 15.2f $ **FLOATING
C5001 li_4468_117244# AVSS 15.2f $ **FLOATING
C5002 li_4468_117404# AVSS 15.2f $ **FLOATING
C5003 li_4468_118204# AVSS 20.2f $ **FLOATING
C5004 a_4308_51566# AVSS 0.491f $ **FLOATING
C5005 a_4308_51918# AVSS 0.389f $ **FLOATING
C5006 xbb1.xa3.M0.D AVSS 0.063f
C5007 xbb1.xa3.M1.D AVSS 0.0143f
C5008 xbb1.xa3.M2.D AVSS 0.0143f
C5009 a_37324_52750# AVSS 0.129f $ **FLOATING
C5010 a_36172_52750# AVSS 0.572f $ **FLOATING
C5011 a_34804_52750# AVSS 0.573f $ **FLOATING
C5012 a_33652_52750# AVSS 0.127f $ **FLOATING
C5013 a_32284_52750# AVSS 0.127f $ **FLOATING
C5014 a_31132_52750# AVSS 0.572f $ **FLOATING
C5015 a_29764_52750# AVSS 0.576f $ **FLOATING
C5016 a_28612_52750# AVSS 0.127f $ **FLOATING
C5017 a_27244_52750# AVSS 0.127f $ **FLOATING
C5018 a_26092_52750# AVSS 0.573f $ **FLOATING
C5019 a_11712_52750# AVSS 0.133f $ **FLOATING
C5020 a_10092_52750# AVSS 0.514f $ **FLOATING
C5021 xbb1.xa3.M3.D AVSS 0.0143f
C5022 a_37324_53102# AVSS 0.00312f $ **FLOATING
C5023 a_36172_53102# AVSS 0.49f $ **FLOATING
C5024 a_34804_53102# AVSS 0.488f $ **FLOATING
C5025 a_33652_53102# AVSS 0.00174f $ **FLOATING
C5026 a_32284_53102# AVSS 0.00174f $ **FLOATING
C5027 a_31132_53102# AVSS 0.49f $ **FLOATING
C5028 a_29764_53102# AVSS 0.488f $ **FLOATING
C5029 a_28612_53102# AVSS 0.00174f $ **FLOATING
C5030 a_27244_53102# AVSS 0.00174f $ **FLOATING
C5031 a_26092_53102# AVSS 0.49f $ **FLOATING
C5032 xbb1.xa3.M4.D AVSS 0.0143f
C5033 xaa4.xa1.M0.D AVSS 0.0804f
C5034 a_37324_53454# AVSS 0.00288f $ **FLOATING
C5035 a_36172_53454# AVSS 0.365f $ **FLOATING
C5036 a_34804_53454# AVSS 0.365f $ **FLOATING
C5037 a_33652_53454# AVSS 0.0015f $ **FLOATING
C5038 a_32284_53454# AVSS 0.0015f $ **FLOATING
C5039 a_31132_53454# AVSS 0.364f $ **FLOATING
C5040 a_29764_53454# AVSS 0.365f $ **FLOATING
C5041 a_28612_53454# AVSS 0.0015f $ **FLOATING
C5042 a_27244_53454# AVSS 0.0015f $ **FLOATING
C5043 a_26092_53454# AVSS 0.365f $ **FLOATING
C5044 xbb1.xa3.M5.D AVSS 0.0143f
C5045 xaa4.xa1.M1.D AVSS 0.0219f
C5046 xaa6.xg.XA1.MN0.D AVSS 0.169f
C5047 xaa6.xf.XA1.MN0.D AVSS 0.169f
C5048 xaa6.xe.XA1.MN0.D AVSS 0.15f
C5049 xaa6.xd.XA1.MN0.D AVSS 0.169f
C5050 xaa6.xc.XA1.MN0.D AVSS 0.15f
C5051 xbb1.xa3.M6.D AVSS 0.0143f
C5052 xaa4.xa1.M2.D AVSS 0.0191f
C5053 a_37324_53806# AVSS 0.00295f $ **FLOATING
C5054 a_36172_53806# AVSS 0.384f $ **FLOATING
C5055 a_34804_53806# AVSS 0.384f $ **FLOATING
C5056 a_33652_53806# AVSS 0.00156f $ **FLOATING
C5057 a_32284_53806# AVSS 0.00156f $ **FLOATING
C5058 a_31132_53806# AVSS 0.383f $ **FLOATING
C5059 a_29764_53806# AVSS 0.384f $ **FLOATING
C5060 a_28612_53806# AVSS 0.00156f $ **FLOATING
C5061 a_27244_53806# AVSS 0.00156f $ **FLOATING
C5062 a_26092_53806# AVSS 0.383f $ **FLOATING
C5063 xbb1.xa3.M7.D AVSS 0.0143f
C5064 xaa4.xa1.M3.D AVSS 0.0178f
C5065 xaa4.xa1.M4.D AVSS 0.0172f
C5066 a_4308_53678# AVSS 0.47f $ **FLOATING
C5067 a_244_52750# AVSS 0.13f $ **FLOATING
C5068 a_n908_52750# AVSS 0.573f $ **FLOATING
C5069 a_244_53102# AVSS 0.00312f $ **FLOATING
C5070 a_n908_53102# AVSS 0.49f $ **FLOATING
C5071 a_244_53454# AVSS 0.00294f $ **FLOATING
C5072 a_n908_53454# AVSS 0.363f $ **FLOATING
C5073 xaa0.xa1.MP1.D AVSS 0.00161f
C5074 a_37324_54158# AVSS 0.00288f $ **FLOATING
C5075 a_36172_54158# AVSS 0.387f $ **FLOATING
C5076 a_34804_54158# AVSS 0.387f $ **FLOATING
C5077 a_33652_54158# AVSS 0.0015f $ **FLOATING
C5078 a_32284_54158# AVSS 0.0015f $ **FLOATING
C5079 a_31132_54158# AVSS 0.387f $ **FLOATING
C5080 a_29764_54158# AVSS 0.387f $ **FLOATING
C5081 a_28612_54158# AVSS 0.0015f $ **FLOATING
C5082 a_27244_54158# AVSS 0.0015f $ **FLOATING
C5083 a_26092_54158# AVSS 0.388f $ **FLOATING
C5084 xaa4.xa1.M5.D AVSS 0.0169f
C5085 xaa4.xa1.M6.D AVSS 0.0166f
C5086 a_11712_54334# AVSS 0.00312f $ **FLOATING
C5087 xaa4.xa1.M7.D AVSS 0.0165f
C5088 a_37324_54510# AVSS 0.00288f $ **FLOATING
C5089 a_36172_54510# AVSS 0.364f $ **FLOATING
C5090 a_34804_54510# AVSS 0.364f $ **FLOATING
C5091 a_33652_54510# AVSS 0.0015f $ **FLOATING
C5092 a_32284_54510# AVSS 0.0015f $ **FLOATING
C5093 a_31132_54510# AVSS 0.364f $ **FLOATING
C5094 a_29764_54510# AVSS 0.364f $ **FLOATING
C5095 a_28612_54510# AVSS 0.0015f $ **FLOATING
C5096 a_27244_54510# AVSS 0.0015f $ **FLOATING
C5097 a_26092_54510# AVSS 0.365f $ **FLOATING
C5098 xaa6.xg.XA3.MP0.D AVSS 0.00886f
C5099 xaa6.xg.XA3.MN0.D AVSS 0.162f
C5100 xaa6.xg.XA3.MN1.G AVSS 1.62f
C5101 xaa6.xf.XA3.MN0.D AVSS 0.162f
C5102 xaa6.xf.XA3.MP0.D AVSS 0.00886f
C5103 xaa6.xe.XA3.MP0.D AVSS 0.00886f
C5104 xaa6.xe.XA3.MN0.D AVSS 0.162f
C5105 xaa6.xd.XA3.MN0.D AVSS 0.162f
C5106 xaa6.xd.XA3.MP0.D AVSS 0.00886f
C5107 xaa6.xc.XA3.MP0.D AVSS 0.00886f
C5108 xaa6.xc.XA3.MN0.D AVSS 0.162f
C5109 a_10092_54510# AVSS 0.372f $ **FLOATING
C5110 a_37324_54862# AVSS 0.00288f $ **FLOATING
C5111 a_36172_54862# AVSS 0.383f $ **FLOATING
C5112 a_34804_54862# AVSS 0.383f $ **FLOATING
C5113 a_33652_54862# AVSS 0.0015f $ **FLOATING
C5114 a_32284_54862# AVSS 0.0015f $ **FLOATING
C5115 a_31132_54862# AVSS 0.383f $ **FLOATING
C5116 a_29764_54862# AVSS 0.383f $ **FLOATING
C5117 a_28612_54862# AVSS 0.0015f $ **FLOATING
C5118 a_27244_54862# AVSS 0.0015f $ **FLOATING
C5119 a_26092_54862# AVSS 0.384f $ **FLOATING
C5120 xaa6.xg.XA4.MN0.G AVSS 0.53f
C5121 a_37324_55214# AVSS 0.00288f $ **FLOATING
C5122 a_36172_55214# AVSS 0.364f $ **FLOATING
C5123 a_34804_55214# AVSS 0.364f $ **FLOATING
C5124 a_33652_55214# AVSS 0.0015f $ **FLOATING
C5125 a_32284_55214# AVSS 0.0015f $ **FLOATING
C5126 a_31132_55214# AVSS 0.364f $ **FLOATING
C5127 a_29764_55214# AVSS 0.364f $ **FLOATING
C5128 a_28612_55214# AVSS 0.0015f $ **FLOATING
C5129 a_27244_55214# AVSS 0.0015f $ **FLOATING
C5130 a_26092_55214# AVSS 0.364f $ **FLOATING
C5131 a_10092_55038# AVSS 0.365f $ **FLOATING
C5132 xaa6.xg.XA4.MP0.D AVSS 0.00592f
C5133 xaa6.xg.XA4.MN0.D AVSS 0.139f
C5134 xaa6.xg.XA4.MP1.G AVSS 0.0255f
C5135 xaa6.xf.XA4.MN0.D AVSS 0.139f
C5136 xaa6.xf.XA4.MP0.D AVSS 0.00592f
C5137 xaa6.xe.XA4.MP0.D AVSS 0.00592f
C5138 xaa6.xe.XA4.MN0.D AVSS 0.139f
C5139 xaa6.xd.XA4.MN0.D AVSS 0.139f
C5140 xaa6.xd.XA4.MP0.D AVSS 0.00592f
C5141 xaa6.xc.XA4.MP0.D AVSS 0.00592f
C5142 xaa6.xc.XA4.MN0.D AVSS 0.139f
C5143 CK_REF AVSS 0.957f
C5144 a_244_53806# AVSS 0.00288f $ **FLOATING
C5145 a_n908_53806# AVSS 0.363f $ **FLOATING
C5146 xaa0.xa1.MN2.D AVSS 0.138f
C5147 xaa0.xa1.MN0.D AVSS 1.16f
C5148 a_244_54158# AVSS 0.00288f $ **FLOATING
C5149 a_n908_54158# AVSS 0.406f $ **FLOATING
C5150 a_244_54510# AVSS 0.00288f $ **FLOATING
C5151 a_n908_54510# AVSS 0.386f $ **FLOATING
C5152 xaa0.xa2a.MN0.G AVSS 1.03f
C5153 a_244_54862# AVSS 0.00288f $ **FLOATING
C5154 a_n908_54862# AVSS 0.384f $ **FLOATING
C5155 a_37324_55566# AVSS 0.00288f $ **FLOATING
C5156 a_36172_55566# AVSS 0.383f $ **FLOATING
C5157 a_34804_55566# AVSS 0.383f $ **FLOATING
C5158 a_33652_55566# AVSS 0.0015f $ **FLOATING
C5159 a_32284_55566# AVSS 0.0015f $ **FLOATING
C5160 a_31132_55566# AVSS 0.383f $ **FLOATING
C5161 a_29764_55566# AVSS 0.383f $ **FLOATING
C5162 a_28612_55566# AVSS 0.0015f $ **FLOATING
C5163 a_27244_55566# AVSS 0.0015f $ **FLOATING
C5164 a_26092_55566# AVSS 0.383f $ **FLOATING
C5165 xaa4.xa1.M8.D AVSS 0.462f
C5166 xaa6.xg.XA5.MN0.G AVSS 1.26f
C5167 xaa6.xg.XA5.MN0.D AVSS 0.229f
C5168 xaa6.xf.XA5.MN0.G AVSS 1.25f
C5169 xaa6.xe.XA5.MN0.G AVSS 1.26f
C5170 xaa6.xd.XA5.MN0.G AVSS 1.25f
C5171 xaa6.xc.XA5.MN0.G AVSS 1.26f
C5172 a_10092_55566# AVSS 0.425f $ **FLOATING
C5173 a_5844_55150# AVSS 0.132f $ **FLOATING
C5174 a_4692_55150# AVSS 0.57f $ **FLOATING
C5175 a_5844_55502# AVSS 0.00337f $ **FLOATING
C5176 a_4692_55502# AVSS 0.49f $ **FLOATING
C5177 xaa4.xa2.M0.D AVSS 0.807f
C5178 a_37324_55918# AVSS 0.00288f $ **FLOATING
C5179 a_36172_55918# AVSS 0.387f $ **FLOATING
C5180 a_34804_55918# AVSS 0.387f $ **FLOATING
C5181 a_33652_55918# AVSS 0.0015f $ **FLOATING
C5182 a_32284_55918# AVSS 0.0015f $ **FLOATING
C5183 a_31132_55918# AVSS 0.387f $ **FLOATING
C5184 a_29764_55918# AVSS 0.387f $ **FLOATING
C5185 a_28612_55918# AVSS 0.0015f $ **FLOATING
C5186 a_27244_55918# AVSS 0.0015f $ **FLOATING
C5187 a_26092_55918# AVSS 0.388f $ **FLOATING
C5188 a_11712_55918# AVSS 0.00667f $ **FLOATING
C5189 xaa6.xg.XA6.MN0.G AVSS 0.523f
C5190 xaa6.xf.XA6.MN0.G AVSS 1.29f
C5191 xaa6.xe.XA6.MN0.G AVSS 1.29f
C5192 xaa6.xd.XA6.MN0.G AVSS 1.29f
C5193 xaa6.xc.XA6.MN0.G AVSS 1.29f
C5194 a_37324_56270# AVSS 0.00288f $ **FLOATING
C5195 a_36172_56270# AVSS 0.362f $ **FLOATING
C5196 a_34804_56270# AVSS 0.362f $ **FLOATING
C5197 a_33652_56270# AVSS 0.0015f $ **FLOATING
C5198 a_32284_56270# AVSS 0.0015f $ **FLOATING
C5199 a_31132_56270# AVSS 0.362f $ **FLOATING
C5200 a_29764_56270# AVSS 0.362f $ **FLOATING
C5201 a_28612_56270# AVSS 0.0015f $ **FLOATING
C5202 a_27244_56270# AVSS 0.0015f $ **FLOATING
C5203 a_26092_56270# AVSS 0.363f $ **FLOATING
C5204 xaa6.xg.XA6.MP0.D AVSS 0.00886f
C5205 xaa6.xg.XA6.MN0.D AVSS 0.146f
C5206 xaa6.xf.XA6.MN0.D AVSS 0.146f
C5207 xaa6.xf.XA6.MP0.D AVSS 0.00886f
C5208 xaa6.xe.XA6.MP0.D AVSS 0.00886f
C5209 xaa6.xe.XA6.MN0.D AVSS 0.146f
C5210 xaa6.xd.XA6.MN0.D AVSS 0.146f
C5211 xaa6.xd.XA6.MP0.D AVSS 0.00886f
C5212 xaa6.xc.XA6.MP0.D AVSS 0.00886f
C5213 xaa6.xc.XA6.MN0.D AVSS 0.146f
C5214 a_5844_55854# AVSS 0.00302f $ **FLOATING
C5215 a_4692_55854# AVSS 0.386f $ **FLOATING
C5216 a_5844_56206# AVSS 0.087f $ **FLOATING
C5217 a_4692_56206# AVSS 0.436f $ **FLOATING
C5218 xaa0.xa1.MN2.S AVSS 1.79f
C5219 a_244_55214# AVSS 0.00288f $ **FLOATING
C5220 a_n908_55214# AVSS 0.367f $ **FLOATING
C5221 xaa0.xa3.MP0.D AVSS 0.00597f
C5222 a_244_55566# AVSS 0.003f $ **FLOATING
C5223 a_n908_55566# AVSS 0.407f $ **FLOATING
C5224 xaa0.xa1.MN0.G AVSS 2.58f
C5225 a_244_55918# AVSS 0.00298f $ **FLOATING
C5226 a_n908_55918# AVSS 0.362f $ **FLOATING
C5227 xaa0.xa5.MP1.D AVSS 0.00161f
C5228 a_37324_56622# AVSS 0.00296f $ **FLOATING
C5229 a_36172_56622# AVSS 0.382f $ **FLOATING
C5230 a_34804_56622# AVSS 0.382f $ **FLOATING
C5231 a_33652_56622# AVSS 0.00158f $ **FLOATING
C5232 a_32284_56622# AVSS 0.00158f $ **FLOATING
C5233 a_31132_56622# AVSS 0.382f $ **FLOATING
C5234 a_29764_56622# AVSS 0.382f $ **FLOATING
C5235 a_28612_56622# AVSS 0.0016f $ **FLOATING
C5236 a_27244_56622# AVSS 0.00158f $ **FLOATING
C5237 a_26092_56622# AVSS 0.382f $ **FLOATING
C5238 a_37324_56974# AVSS 0.00286f $ **FLOATING
C5239 a_36172_56974# AVSS 0.362f $ **FLOATING
C5240 a_34804_56974# AVSS 0.362f $ **FLOATING
C5241 a_33652_56974# AVSS 0.00147f $ **FLOATING
C5242 a_32284_56974# AVSS 0.00147f $ **FLOATING
C5243 a_31132_56974# AVSS 0.362f $ **FLOATING
C5244 a_29764_56974# AVSS 0.362f $ **FLOATING
C5245 a_28612_56974# AVSS 0.00151f $ **FLOATING
C5246 a_27244_56974# AVSS 0.00147f $ **FLOATING
C5247 a_26092_56974# AVSS 0.363f $ **FLOATING
C5248 xaa6.xg.XA7.MN2.D AVSS 0.181f
C5249 xaa6.xg.XA7.MN0.G AVSS 0.51f
C5250 xaa6.xf.XA7.MN2.D AVSS 0.181f
C5251 xaa6.xe.XA7.MN2.D AVSS 0.181f
C5252 xaa6.xd.XA7.MN2.D AVSS 0.181f
C5253 xaa6.xc.XA7.MN2.D AVSS 0.181f
C5254 a_244_56270# AVSS 0.00307f $ **FLOATING
C5255 a_n908_56270# AVSS 0.362f $ **FLOATING
C5256 xaa0.xa5.MN2.D AVSS 0.152f
C5257 xaa0.xa5.MN0.D AVSS 1.16f
C5258 a_244_56622# AVSS 0.00348f $ **FLOATING
C5259 a_n908_56622# AVSS 0.407f $ **FLOATING
C5260 xaa0.xa3.MN1.G AVSS 2.02f
C5261 a_244_56974# AVSS 0.129f $ **FLOATING
C5262 a_n908_56974# AVSS 0.465f $ **FLOATING
C5263 a_37324_57326# AVSS 0.00293f $ **FLOATING
C5264 a_36172_57326# AVSS 0.359f $ **FLOATING
C5265 a_34804_57326# AVSS 0.359f $ **FLOATING
C5266 a_33652_57326# AVSS 0.00155f $ **FLOATING
C5267 a_32284_57326# AVSS 0.00155f $ **FLOATING
C5268 a_31132_57326# AVSS 0.359f $ **FLOATING
C5269 a_29764_57326# AVSS 0.359f $ **FLOATING
C5270 a_28612_57326# AVSS 0.00162f $ **FLOATING
C5271 a_27244_57326# AVSS 0.00155f $ **FLOATING
C5272 a_26092_57326# AVSS 0.36f $ **FLOATING
C5273 xaa6.xg.XA7.MN0.D AVSS 0.248f
C5274 xaa6.xg.XA7.MP1.G AVSS 1.85f
C5275 xaa6.xg.XA7.MN1.G AVSS 1.35f
C5276 xaa6.xf.XA7.MN0.D AVSS 0.248f
C5277 xaa6.xf.XA7.MN1.G AVSS 2.9f
C5278 xaa6.xf.XA7.MP1.G AVSS 1.85f
C5279 xaa6.xe.XA7.MN0.D AVSS 0.248f
C5280 xaa6.xe.XA7.MP1.G AVSS 1.85f
C5281 xaa6.xe.XA7.MN1.G AVSS 2.91f
C5282 xaa6.xd.XA7.MN0.D AVSS 0.248f
C5283 xaa6.xd.XA7.MN1.G AVSS 2.9f
C5284 xaa6.xd.XA7.MP1.G AVSS 1.85f
C5285 xaa6.xc.XA7.MN0.D AVSS 0.248f
C5286 xaa6.xc.XA7.MP1.G AVSS 1.85f
C5287 xaa6.xc.XA7.MN1.G AVSS 3.02f
C5288 a_11712_57502# AVSS 0.00378f $ **FLOATING
C5289 a_37324_57678# AVSS 0.00341f $ **FLOATING
C5290 a_36172_57678# AVSS 0.381f $ **FLOATING
C5291 a_34804_57678# AVSS 0.381f $ **FLOATING
C5292 a_33652_57678# AVSS 0.00203f $ **FLOATING
C5293 a_32284_57678# AVSS 0.00203f $ **FLOATING
C5294 a_31132_57678# AVSS 0.381f $ **FLOATING
C5295 a_29764_57678# AVSS 0.381f $ **FLOATING
C5296 a_28612_57678# AVSS 0.00222f $ **FLOATING
C5297 a_27244_57678# AVSS 0.00203f $ **FLOATING
C5298 a_26092_57678# AVSS 0.382f $ **FLOATING
C5299 xaa6.xg.XA7.MN1.D AVSS 2.68f
C5300 xaa6.xf.XA1.MN0.G AVSS 2.93f
C5301 xaa6.xf.XA7.MN1.D AVSS 2.67f
C5302 xaa6.xe.XA1.MN0.G AVSS 2.89f
C5303 xaa6.xe.XA7.MN1.D AVSS 2.68f
C5304 xaa6.xd.XA1.MN0.G AVSS 3.54f
C5305 xaa6.xd.XA7.MN1.D AVSS 2.67f
C5306 xaa6.xc.XA1.MN0.G AVSS 3.02f
C5307 xaa6.xc.XA7.MN1.D AVSS 2.67f
C5308 xaa0.xa5.MN2.G AVSS 15.4f
C5309 a_37324_58030# AVSS 0.129f $ **FLOATING
C5310 a_36172_58030# AVSS 0.462f $ **FLOATING
C5311 a_34804_58030# AVSS 0.463f $ **FLOATING
C5312 a_33652_58030# AVSS 0.127f $ **FLOATING
C5313 a_32284_58030# AVSS 0.127f $ **FLOATING
C5314 a_31132_58030# AVSS 0.462f $ **FLOATING
C5315 a_29764_58030# AVSS 0.463f $ **FLOATING
C5316 a_28612_58030# AVSS 0.131f $ **FLOATING
C5317 a_27244_58030# AVSS 0.127f $ **FLOATING
C5318 a_26092_58030# AVSS 0.465f $ **FLOATING
C5319 a_5844_57790# AVSS 0.109f $ **FLOATING
C5320 a_4692_57790# AVSS 0.472f $ **FLOATING
C5321 xaa3.xa1capd.B AVSS 5.24f
C5322 a_5844_58142# AVSS 0.00346f $ **FLOATING
C5323 a_4692_58142# AVSS 0.385f $ **FLOATING
C5324 xaa3.xa2.MN0.D AVSS 1.17f
C5325 a_5844_58494# AVSS 0.0871f $ **FLOATING
C5326 a_4692_58494# AVSS 0.436f $ **FLOATING
C5327 a_11712_59086# AVSS 0.00667f $ **FLOATING
C5328 a_640_59750# AVSS 0.13f $ **FLOATING
C5329 a_n908_59750# AVSS 0.519f $ **FLOATING
C5330 xaa4.xa4.M0.D AVSS 1.41f
C5331 a_11712_60670# AVSS 0.0913f $ **FLOATING
C5332 a_29764_60750# AVSS 0.493f $ **FLOATING
C5333 a_28612_60750# AVSS 0.136f $ **FLOATING
C5334 a_27244_60750# AVSS 0.127f $ **FLOATING
C5335 a_26092_60750# AVSS 0.492f $ **FLOATING
C5336 a_5844_60078# AVSS 0.109f $ **FLOATING
C5337 a_4692_60078# AVSS 0.472f $ **FLOATING
C5338 xaa1.xb1.M0.D AVSS 1.41e-25
C5339 xaa3.xa3a.MN0.D AVSS 5.25f
C5340 xaa1.xa1.M0.D AVSS 0.0851f
C5341 a_640_60278# AVSS 0.00372f $ **FLOATING
C5342 xaa1.xa1.M1.D AVSS 0.0262f
C5343 a_5844_60430# AVSS 0.00346f $ **FLOATING
C5344 a_4692_60430# AVSS 0.385f $ **FLOATING
C5345 xaa3.xa4.MN0.D AVSS 1.17f
C5346 xaa1.xa1.M2.D AVSS 0.0234f
C5347 xaa1.xb2.M0.D AVSS 2.93e-25
C5348 a_5844_60782# AVSS 0.0871f $ **FLOATING
C5349 a_4692_60782# AVSS 0.436f $ **FLOATING
C5350 xaa1.xa1.M3.D AVSS 0.0222f
C5351 a_640_60806# AVSS 0.00352f $ **FLOATING
C5352 xaa1.xa1.M4.D AVSS 0.0216f
C5353 xaa1.xb2.M7.D AVSS 1.28e-24
C5354 a_29764_61102# AVSS 0.366f $ **FLOATING
C5355 a_28612_61102# AVSS 0.00226f $ **FLOATING
C5356 a_27244_61102# AVSS 0.00182f $ **FLOATING
C5357 a_26092_61102# AVSS 0.384f $ **FLOATING
C5358 xaa0.xa2a.MN0.D AVSS 3.65f
C5359 xaa1.xa1.M5.D AVSS 0.0212f
C5360 xaa5.xb1.MN0.D AVSS 0.175f
C5361 xaa5.xa3.xc1a.D AVSS 0.00756f
C5362 a_640_61158# AVSS 0.00348f $ **FLOATING
C5363 xaa1.xa1.M6.D AVSS 0.021f
C5364 a_29764_61454# AVSS 0.38f $ **FLOATING
C5365 a_28612_61454# AVSS 0.00177f $ **FLOATING
C5366 a_27244_61454# AVSS 0.00161f $ **FLOATING
C5367 a_26092_61454# AVSS 0.389f $ **FLOATING
C5368 PWRUP_1V8 AVSS 37f
C5369 xaa1.xa1.M7.D AVSS 0.0209f
C5370 xaa1.xa1.M8.D AVSS 0.735f
C5371 xaa5.xb1.MN1.D AVSS 0.983f
C5372 a_640_61510# AVSS 0.092f $ **FLOATING
C5373 a_n908_61510# AVSS 0.398f $ **FLOATING
C5374 a_29764_61806# AVSS 0.384f $ **FLOATING
C5375 a_28612_61806# AVSS 0.00163f $ **FLOATING
C5376 a_27244_61806# AVSS 0.00152f $ **FLOATING
C5377 a_26092_61806# AVSS 0.388f $ **FLOATING
C5378 xaa1.xa2.M0.D AVSS 0.0691f
C5379 xaa5.xb2_0.MN0.D AVSS 0.897f
C5380 xaa5.xa3.xc2a.D AVSS 0.00756f
C5381 xaa1.xa2.M1.D AVSS 0.0204f
C5382 a_29764_62158# AVSS 0.384f $ **FLOATING
C5383 a_28612_62158# AVSS 0.00158f $ **FLOATING
C5384 a_27244_62158# AVSS 0.00151f $ **FLOATING
C5385 a_26092_62158# AVSS 0.384f $ **FLOATING
C5386 xaa1.xa2.M2.D AVSS 0.0204f
C5387 xaa5.xb2_1.MN0.D AVSS 0.893f
C5388 xaa5.xa3.xb1_0.D AVSS 1.91f
C5389 xaa5.xa4.MN0.D AVSS 0.216f
C5390 a_29764_62510# AVSS 0.384f $ **FLOATING
C5391 a_28612_62510# AVSS 0.00149f $ **FLOATING
C5392 a_27244_62510# AVSS 0.00152f $ **FLOATING
C5393 a_26092_62510# AVSS 0.388f $ **FLOATING
C5394 xaa5.xb2_2.MN0.D AVSS 0.893f
C5395 xaa5.xa3.xb2_0.D AVSS 1.43f
C5396 CK AVSS 13.3f
C5397 a_29764_62862# AVSS 0.384f $ **FLOATING
C5398 a_28612_62862# AVSS 0.00149f $ **FLOATING
C5399 a_27244_62862# AVSS 0.00159f $ **FLOATING
C5400 a_26092_62862# AVSS 0.467f $ **FLOATING
C5401 xaa5.xb2_3.MN0.D AVSS 0.893f
C5402 a_29764_63214# AVSS 0.384f $ **FLOATING
C5403 a_28612_63214# AVSS 0.00149f $ **FLOATING
C5404 a_27244_63214# AVSS 0.0893f $ **FLOATING
C5405 a_26092_63214# AVSS 0.531f $ **FLOATING
C5406 a_5844_62366# AVSS 0.109f $ **FLOATING
C5407 a_4692_62366# AVSS 0.472f $ **FLOATING
C5408 xaa1.xa2.M3.D AVSS 0.0204f
C5409 xaa3.xa5a.MN0.D AVSS 5.25f
C5410 xaa1.xa2.M4.D AVSS 0.0204f
C5411 a_5844_62718# AVSS 0.00352f $ **FLOATING
C5412 a_4692_62718# AVSS 0.385f $ **FLOATING
C5413 xaa1.xa2.M5.D AVSS 0.0204f
C5414 xaa3.xa6.MN0.D AVSS 1.11f
C5415 xaa1.xa2.M6.D AVSS 0.0204f
C5416 a_5844_63070# AVSS 0.00312f $ **FLOATING
C5417 a_4692_63070# AVSS 0.384f $ **FLOATING
C5418 xaa1.xa2.M7.D AVSS 0.0204f
C5419 xaa5.xb2_4.MN0.D AVSS 0.893f
C5420 a_29764_63566# AVSS 0.381f $ **FLOATING
C5421 a_28612_63566# AVSS 0.00266f $ **FLOATING
C5422 xaa5.xa3.xb2_0.G AVSS 3.22f
C5423 a_29764_63918# AVSS 0.381f $ **FLOATING
C5424 a_28612_63918# AVSS 0.00266f $ **FLOATING
C5425 xaa4.xa2.M0.G AVSS 0.791p
C5426 xaa5.xa3.xb1_0.G AVSS 3.71f
C5427 xaa5.xb1.MN1.G AVSS 2.59f
C5428 xaa3.xa1b.MN0.D AVSS 7.1f
C5429 IBPSR_1U AVSS 23.7f
C5430 a_n908_63270# AVSS 0.367f $ **FLOATING
C5431 a_5844_63422# AVSS 0.00312f $ **FLOATING
C5432 a_4692_63422# AVSS 0.369f $ **FLOATING
C5433 xaa1.xa2.M8.D AVSS 0.166f
C5434 xaa3.xa8.MP0.D AVSS 0.00592f
C5435 xaa3.xa7.MN0.D AVSS 1.03f
C5436 xaa0.xa6.MN0.D AVSS 3.79f
C5437 a_n908_63622# AVSS 0.384f $ **FLOATING
C5438 a_5844_63774# AVSS 0.00349f $ **FLOATING
C5439 a_4692_63774# AVSS 0.407f $ **FLOATING
C5440 xaa3.xa9.MN0.D AVSS 0.29f
C5441 a_5844_64126# AVSS 0.129f $ **FLOATING
C5442 a_4692_64126# AVSS 0.468f $ **FLOATING
C5443 xaa1.xa4.M0.G AVSS 5.85f
C5444 a_n908_64150# AVSS 0.487f $ **FLOATING
C5445 a_29764_64270# AVSS 0.469f $ **FLOATING
C5446 a_28612_64270# AVSS 0.00291f $ **FLOATING
C5447 xaa5.xb3.MP1.D AVSS 0.119f
C5448 a_29764_64622# AVSS 0.568f $ **FLOATING
C5449 a_28612_64622# AVSS 0.128f $ **FLOATING
C5450 a_2948_70022# AVSS 2.59f $ **FLOATING
C5451 xaa1.xa3.D AVSS 0.309p
C5452 a_2084_70022# AVSS 0.843f
C5453 a_1652_72222# AVSS 1.08f
C5454 a_1220_70022# AVSS 0.778f
C5455 a_788_72222# AVSS 1.08f
C5456 a_356_70022# AVSS 0.778f
C5457 a_n76_72222# AVSS 1.08f
C5458 a_n508_70022# AVSS 0.843f
C5459 a_n940_70022# AVSS 2.59f $ **FLOATING
C5460 a_2948_74698# AVSS 2.59f $ **FLOATING
C5461 xaa1.xa4.M0.D AVSS 4.98p
C5462 a_2084_74698# AVSS 0.843f
C5463 a_1652_76898# AVSS 1.08f
C5464 a_1220_74698# AVSS 0.778f
C5465 a_788_76898# AVSS 1.08f
C5466 a_356_74698# AVSS 0.778f
C5467 a_n76_76898# AVSS 1.08f
C5468 a_n508_74698# AVSS 0.843f
C5469 xbb0.xa1.XA1.N AVSS 3.4f
C5470 a_n940_74698# AVSS 2.59f $ **FLOATING
C5471 AVDD AVSS 0.418p
.ends

