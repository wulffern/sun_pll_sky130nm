** sch_path: /Users/wulff/pro/aicex/ip/sun_pll_sky130nm/work/../design/SUN_PLL_SKY130NM/SUN_PLL.sch
.subckt SUN_PLL AVDD AVSS PWRUP_1V8 CK_REF CK IBPSR_1U
*.ipin AVDD
*.ipin AVSS
*.ipin PWRUP_1V8
*.ipin CK_REF
*.opin CK
*.ipin IBPSR_1U
xa0 AVDD CP_UP_N CK_REF CP_DOWN CK_FB AVSS SUN_PLL_PFD
xa1 AVDD CP_UP_N VLPF CP_DOWN IBPSR_1U AVSS VLPFZ PWRUP_1V8 KICK SUN_PLL_CP
xa4 AVDD VDD_ROSC VLPF VDD_ROSC IBPSR_1U AVSS SUN_PLL_BUF
xa5 AVDD CK VDD_ROSC PWRUP_1V8 AVSS SUN_PLL_ROSC
xaa3 AVDD KICK net1 PWRUP_1V8 AVSS PWRUP_1V8_N SUN_PLL_KICK
xaa6 AVDD CK_FB CK PWRUP_1V8 AVSS SUN_PLL_DIVN
xbb1 IBPSR_1U PWRUP_1V8_N AVSS SUN_PLL_BIAS
xd0 VLPFZ AVSS VLPF SUN_PLL_LPF
.ends

* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_ROSC.sym # of pins=5
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_ROSC.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_ROSC.sch
.subckt SUN_PLL_ROSC AVDD CK VDD_ROSC PWRUP_1V8 AVSS
*.ipin AVDD
*.opin CK
*.ipin VDD_ROSC
*.ipin PWRUP_1V8
*.ipin AVSS
xa3 N_2 N_1 CKUP CKDWN AVDD AVSS SUN_PLL_LSCORE
xa4 CKDWN NC1 AVDD AVSS SUNTR_IVX1_CV
xa5 CKUP CK AVDD AVSS SUNTR_IVX1_CV
xa6 AVDD AVSS SUNTR_TAPCELLB_CV
xb1 PWRUP_1V8 N_0 NI AVDD AVSS VDD_ROSC AVSS SUNTRB_NDX1_CV
xb2_0 NI N_7 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_1 N_7 N_6 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_2 N_6 N_5 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_3 N_5 N_4 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_4 N_4 N_3 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_5 N_3 N_2 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_6 N_2 N_1 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb2_7 N_1 N_0 AVDD AVSS VDD_ROSC AVSS SUNTRB_IVX1_CV
xb3 AVDD AVSS SUNTRB_TAPCELLBAVSS_CV
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_DIVN.sym # of pins=5
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_DIVN.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_DIVN.sch
.subckt SUN_PLL_DIVN AVDD CK_FB CK PWRUP_1V8 AVSS
*.ipin PWRUP_1V8
*.ipin CK
*.ipin AVDD
*.ipin AVSS
*.opin CK_FB
xc N2 D2 PWRUP_1V8 CK_FB N2 AVDD AVSS SUNTR_DFRNQNX1_CV
xd N3 D3 PWRUP_1V8 D2 N3 AVDD AVSS SUNTR_DFRNQNX1_CV
xe N4 D4 PWRUP_1V8 D3 N4 AVDD AVSS SUNTR_DFRNQNX1_CV
xf N5 D5 PWRUP_1V8 D4 N5 AVDD AVSS SUNTR_DFRNQNX1_CV
xg N6 CK PWRUP_1V8 D5 N6 AVDD AVSS SUNTR_DFRNQNX1_CV
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_BIAS.sym # of pins=3
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_BIAS.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_BIAS.sch
.subckt SUN_PLL_BIAS IBPSR_1U PWRUP_1V8_N AVSS
*.ipin IBPSR_1U
*.ipin PWRUP_1V8_N
*.ipin AVSS
xa2 IBPSR_1U PWRUP_1V8_N AVSS AVSS SUNTR_NCHDL
xa3 IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_BUF.sym # of pins=6
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_BUF.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_BUF.sch
.subckt SUN_PLL_BUF AVDD VFB VI VO VBN AVSS
*.ipin AVDD
*.ipin VFB
*.ipin VI
*.opin VO
*.ipin VBN
*.ipin AVSS
xa1 VS VBN AVSS AVSS SUNTR_NCHDLCM
xa2 VDP VFB VS AVSS SUNTR_NCHDLA
xa4 VGP VI VS AVSS SUNTR_NCHDLA
xc1_0 VGP VDP AVDD AVDD SUNTR_PCHL
xc1_1 VGP VDP AVDD AVDD SUNTR_PCHL
xc1_2 VGP VDP AVDD AVDD SUNTR_PCHL
xc1_3 VGP VDP AVDD AVDD SUNTR_PCHL
xc2_0 VDP VDP AVDD AVDD SUNTR_PCHL
xc2_1 VDP VDP AVDD AVDD SUNTR_PCHL
xc2_2 VDP VDP AVDD AVDD SUNTR_PCHL
xc2_3 VDP VDP AVDD AVDD SUNTR_PCHL
xc3_0 VO VGP AVDD AVDD SUNTR_PCHL
xc3_1 VO VGP AVDD AVDD SUNTR_PCHL
xc3_10 VO VGP AVDD AVDD SUNTR_PCHL
xc3_2 VO VGP AVDD AVDD SUNTR_PCHL
xc3_3 VO VGP AVDD AVDD SUNTR_PCHL
xc3_4 VO VGP AVDD AVDD SUNTR_PCHL
xc3_5 VO VGP AVDD AVDD SUNTR_PCHL
xc3_6 VO VGP AVDD AVDD SUNTR_PCHL
xc3_7 VO VGP AVDD AVDD SUNTR_PCHL
xc3_8 VO VGP AVDD AVDD SUNTR_PCHL
xc3_9 VO VGP AVDD AVDD SUNTR_PCHL
xd2 VO AVSS SUNSAR_CAP_BSSW_CV
xd3_0 VO AVSS SUNSAR_CAP_BSSW_CV
xd3_1 VO AVSS SUNSAR_CAP_BSSW_CV
xd3_2 VO AVSS SUNSAR_CAP_BSSW_CV
xd3_3 VO AVSS SUNSAR_CAP_BSSW_CV
xd3_4 VO AVSS SUNSAR_CAP_BSSW_CV
xd3_5 VO AVSS SUNSAR_CAP_BSSW_CV
xd3_6 VO AVSS SUNSAR_CAP_BSSW_CV
xd3_7 VO AVSS SUNSAR_CAP_BSSW_CV
xd3_8 VO AVSS SUNSAR_CAP_BSSW_CV
xd3_9 VO AVSS SUNSAR_CAP_BSSW_CV
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_LPF.sym # of pins=3
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_LPF.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_LPF.sch
.subckt SUN_PLL_LPF VLPFZ AVSS VLPF
*.ipin VLPF
*.ipin AVSS
*.ipin VLPFZ
xa1 VN5 VLPF AVSS SUNTR_RPPO8
xa2 VN5 VLPFZ AVSS SUNTR_RPPO8
xb1 VLPF AVSS CAP_LPF
xb2_0 VLPF AVSS CAP_LPF
xb2_1 VLPF AVSS CAP_LPF
xb3_0 VLPFZ AVSS CAP_LPF
xb3_1 VLPFZ AVSS CAP_LPF
xb3_10 VLPFZ AVSS CAP_LPF
xb3_11 VLPFZ AVSS CAP_LPF
xb3_12 VLPFZ AVSS CAP_LPF
xb3_13 VLPFZ AVSS CAP_LPF
xb3_14 VLPFZ AVSS CAP_LPF
xb3_15 VLPFZ AVSS CAP_LPF
xb3_16 VLPFZ AVSS CAP_LPF
xb3_17 VLPFZ AVSS CAP_LPF
xb3_18 VLPFZ AVSS CAP_LPF
xb3_19 VLPFZ AVSS CAP_LPF
xb3_2 VLPFZ AVSS CAP_LPF
xb3_20 VLPFZ AVSS CAP_LPF
xb3_21 VLPFZ AVSS CAP_LPF
xb3_3 VLPFZ AVSS CAP_LPF
xb3_4 VLPFZ AVSS CAP_LPF
xb3_5 VLPFZ AVSS CAP_LPF
xb3_6 VLPFZ AVSS CAP_LPF
xb3_7 VLPFZ AVSS CAP_LPF
xb3_8 VLPFZ AVSS CAP_LPF
xb3_9 VLPFZ AVSS CAP_LPF
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_CP.sym # of pins=9
** sym_path: /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_CP.sym
** sch_path: /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_CP.sch
.subckt SUN_PLL_CP AVDD CP_UP_N LPF CP_DOWN VBN AVSS LPFZ PWRUP_1V8 KICK
*.ipin AVDD
*.ipin CP_UP_N
*.ipin CP_DOWN
*.ipin VBN
*.ipin AVSS
*.opin LPF
*.ipin PWRUP_1V8
*.opin LPFZ
*.ipin KICK
xa1 VBP VBN AVSS AVSS SUNTR_NCHDLCM
xa2 VNS VBN AVSS AVSS SUNTR_NCHDLCM
xa3 LPF CP_DOWN VNS AVSS SUNTR_NCHDL
xa4 LPFZ KICK AVSS AVSS SUNTR_NCHDLA
xb1 VBP VBP AVDD AVDD SUNTR_PCHDLCM
xb2 VPS VBP AVDD AVDD SUNTR_PCHDLCM
xb3 LPF CP_UP_N VPS AVDD SUNTR_PCHDL
xb4 LPF PWRUP_1V8 AVDD AVDD SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_PFD.sym # of pins=6
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_PFD.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_PFD.sch
.subckt SUN_PLL_PFD AVDD CP_UP_N CK_REF CP_DOWN CK_FB AVSS
*.ipin AVDD
*.opin CP_UP_N
*.ipin CK_REF
*.opin CP_DOWN
*.ipin CK_FB
*.ipin AVSS
xa0 AVDD AVSS SUNTR_TAPCELLB_CV
xa1 CFB CK_REF CP_DUP_N AVDD AVSS SUNTR_DFTSPCX1_CV
xa2 CP_DUP_N CP_UP AVDD AVSS SUNTR_IVX1_CV
xa2a CP_UP CP_UP_N AVDD AVSS SUNTR_IVX1_CV
xa3 CP_DUP_N CP_DOWN_N CFB AVDD AVSS SUNTR_NRX1_CV
xa5 CFB CK_FB CP_DOWN_N AVDD AVSS SUNTR_DFTSPCX1_CV
xa6 CP_DOWN_N CP_DOWN AVDD AVSS SUNTR_IVX1_CV
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_KICK.sym # of pins=6
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_KICK.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_KICK.sch
.subckt SUN_PLL_KICK AVDD KICK KICK_N PWRUP_1V8 AVSS PWRUP_1V8_N
*.ipin PWRUP_1V8
*.opin KICK
*.opin KICK_N
*.ipin AVDD
*.ipin AVSS
*.opin PWRUP_1V8_N
xa1a AVDD AVSS SUNTR_TAPCELLB_CV
xa1b PWRUP_1V8 PWRUP_1V8_N AVDD AVSS SUNTR_IVX1_CV
xa1c PWRUP_1V8_N N1 AVDD AVSS SUNTR_IVX1_CV
xa2 N1 N4 AVDD AVSS SUNTR_IVX1_CV
xa5a N4 N5 AVDD AVSS SUNTR_IVX1_CV
xa5capb AVSS N5 SUNTR_DCAPX1_CV
xa6 N5 N6 AVDD AVSS SUNTR_IVX1_CV
xa7 N6 N7 AVDD AVSS SUNTR_IVX1_CV
xa8 PWRUP_1V8_N N7 KICK AVDD AVSS SUNTR_NRX1_CV
xa9 KICK KICK_N AVDD AVSS SUNTR_IVX1_CV
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_IVX1_CV.sym # of pins=4
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV.sch
.subckt SUNTR_IVX1_CV A Y AVDD AVSS
*.ipin A
*.opin Y
*.ipin AVDD
*.ipin AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/SUN_PLL_LSCORE.sym # of pins=6
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_LSCORE.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/SUN_PLL_LSCORE.sch
.subckt SUN_PLL_LSCORE A AN YN Y AVDD AVSS
*.ipin AVDD
*.ipin A
*.ipin AN
*.opin Y
*.opin YN
*.ipin AVSS
xb1_0 Y AN AVSS AVSS SUNTR_NCHDL
xb1_1 Y AN AVSS AVSS SUNTR_NCHDL
xb2_0 YN A AVSS AVSS SUNTR_NCHDL
xb2_1 YN A AVSS AVSS SUNTR_NCHDL
xc1a net2 YN AVDD AVDD SUNTR_PCHDL
xc1b Y YN net2 AVDD SUNTR_PCHDL
xc2a net1 Y AVDD AVDD SUNTR_PCHDL
xc2b YN Y net1 AVDD SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_TAPCELLB_CV.sym # of pins=2
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_TAPCELLB_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_TAPCELLB_CV.sch
.subckt SUNTR_TAPCELLB_CV AVDD AVSS
*.iopin AVDD
*.iopin AVSS
XMN1 AVSS AVSS AVSS AVSS SUNTR_NCHDL
XMP1 AVDD AVDD AVDD AVDD SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_TRB_SKY130NM/SUNTRB_IVX1_CV.sym # of pins=6
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_trb_sky130nm/design/SUN_TRB_SKY130NM/SUNTRB_IVX1_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_trb_sky130nm/design/SUN_TRB_SKY130NM/SUNTRB_IVX1_CV.sch
.subckt SUNTRB_IVX1_CV A Y BULKP BULKN AVDD AVSS
*.ipin A
*.opin Y
*.ipin BULKP
*.ipin BULKN
*.ipin AVDD
*.ipin AVSS
XMN0 Y A AVSS BULKN SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNTRB_PCHDL
.ends


* expanding   symbol:  SUN_TRB_SKY130NM/SUNTRB_NDX1_CV.sym # of pins=7
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_trb_sky130nm/design/SUN_TRB_SKY130NM/SUNTRB_NDX1_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_trb_sky130nm/design/SUN_TRB_SKY130NM/SUNTRB_NDX1_CV.sch
.subckt SUNTRB_NDX1_CV A B Y BULKP BULKN AVDD AVSS
*.ipin A
*.ipin B
*.opin Y
*.ipin BULKP
*.ipin BULKN
*.ipin AVDD
*.ipin AVSS
XMN0 N1 A AVSS BULKN SUNTRB_NCHDL
XMN1 Y B N1 BULKN SUNTRB_NCHDL
XMP0 Y A AVDD BULKP SUNTRB_PCHDL
XMP1 AVDD B Y BULKP SUNTRB_PCHDL
.ends


* expanding   symbol:  SUN_TRB_SKY130NM/SUNTRB_TAPCELLBAVSS_CV.sym # of pins=2
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_trb_sky130nm/design/SUN_TRB_SKY130NM/SUNTRB_TAPCELLBAVSS_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_trb_sky130nm/design/SUN_TRB_SKY130NM/SUNTRB_TAPCELLBAVSS_CV.sch
.subckt SUNTRB_TAPCELLBAVSS_CV AVDD AVSS
*.iopin AVDD
*.iopin AVSS
XMN1 AVSS AVSS AVSS AVSS SUNTRB_NCHDL
XMP1 NC1 NC1 NC1 AVDD SUNTRB_PCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV.sym # of pins=7
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV.sch
.subckt SUNTR_DFRNQNX1_CV D CK RN Q QN AVDD AVSS
*.iopin D
*.iopin CK
*.iopin RN
*.iopin Q
*.iopin QN
*.iopin AVDD
*.iopin AVSS
XXA0 AVDD AVSS SUNTR_TAPCELLB_CV
XXA1 CK RN CKN AVDD AVSS SUNTR_NDX1_CV
XXA2 CKN CKB AVDD AVSS SUNTR_IVX1_CV
XXA3 D CKN CKB A0 AVDD AVSS SUNTR_IVTRIX1_CV
XXA4 A1 CKB CKN A0 AVDD AVSS SUNTR_IVTRIX1_CV
XXA5 A0 A1 AVDD AVSS SUNTR_IVX1_CV
XXA6 A1 CKB CKN QN AVDD AVSS SUNTR_IVTRIX1_CV
XXA7 Q CKN CKB RN QN AVDD AVSS SUNTR_NDTRIX1_CV
XXA8 QN Q AVDD AVSS SUNTR_IVX1_CV
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NCHDLCM.sym # of pins=4
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM.sch
.subckt SUNTR_NCHDLCM D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM0 N0 G S B SUNTR_NCHDL
XM1 N1 G N0 B SUNTR_NCHDL
XM2 N2 G N1 B SUNTR_NCHDL
XM3 N3 G N2 B SUNTR_NCHDL
XM4 N4 G N3 B SUNTR_NCHDL
XM5 N5 G N4 B SUNTR_NCHDL
XM6 N6 G N5 B SUNTR_NCHDL
XM7 N7 G N6 B SUNTR_NCHDL
XM8 D G N7 B SUNTR_NCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NCHDL.sym # of pins=4
** sym_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL.sym
** sch_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL.sch
.subckt SUNTR_NCHDL D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.18 W=1.08 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'  sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NCHDLA.sym # of pins=4
** sym_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA.sym
** sch_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA.sch
.subckt SUNTR_NCHDLA D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM0 D G S B SUNTR_NCHDL
XM1 S G D B SUNTR_NCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_PCHL.sym # of pins=4
** sym_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHL.sym
** sch_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHL.sch
.subckt SUNTR_PCHL D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.36 W=1.08 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'  sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV.sym # of pins=2
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_sar9b_sky130nm/design/SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV.sch
.subckt SUNSAR_CAP_BSSW_CV A B
*.iopin A
*.iopin B
R1 A NC0 sky130_fd_pr__res_generic_m3 W=0.44 L=0.36 m=1
R2 B NC1 sky130_fd_pr__res_generic_m3 W=0.44 L=0.36 m=1
.ends


* expanding   symbol:  SUN_PLL_SKY130NM/CAP_LPF.sym # of pins=2
** sym_path: /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/CAP_LPF.sym
** sch_path: /Users/wulff/data/2023/aicex/ip/sun_pll_sky130nm/design/SUN_PLL_SKY130NM/CAP_LPF.sch
.subckt CAP_LPF A B
*.iopin A
*.iopin B
R1 A NC0 sky130_fd_pr__res_generic_m3 W=0.4 L=0.4 m=1
R2 B NC1 sky130_fd_pr__res_generic_m3 W=0.4 L=0.4 m=1
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_RPPO8.sym # of pins=3
** sym_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8.sym
** sch_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8.sch
.subckt SUNTR_RPPO8 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B SUNTR_RES8
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_PCHDLCM.sym # of pins=4
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLCM.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLCM.sch
.subckt SUNTR_PCHDLCM D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM0 N0 G S B SUNTR_PCHDL
XM7 D G N0 B SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_PCHDL.sym # of pins=4
** sym_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL.sym
** sch_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL.sch
.subckt SUNTR_PCHDL D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.18 W=1.08 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'  sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NRX1_CV.sym # of pins=5
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NRX1_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NRX1_CV.sch
.subckt SUNTR_NRX1_CV A B Y AVDD AVSS
*.iopin A
*.iopin B
*.iopin Y
*.iopin AVDD
*.iopin AVSS
XMN0 Y A AVSS AVSS SUNTR_NCHDL
XMN1 AVSS B Y AVSS SUNTR_NCHDL
XMP0 N1 A AVDD AVDD SUNTR_PCHDL
XMP1 Y B N1 AVDD SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_DFTSPCX1_CV.sym # of pins=5
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFTSPCX1_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFTSPCX1_CV.sch
.subckt SUNTR_DFTSPCX1_CV D CK Q AVDD AVSS
*.iopin D
*.iopin CK
*.iopin Q
*.iopin AVDD
*.iopin AVSS
XMN0 N1 D AVSS AVSS SUNTR_NCHDL
XMN1 AVSS N1 N2 AVSS SUNTR_NCHDL
XMN2 N2 CK Q AVSS SUNTR_NCHDL
XMP0 N1 CK N3 AVDD SUNTR_PCHDL
XMP1 N3 D AVDD AVDD SUNTR_PCHDL
XMP2 Q N1 AVDD AVDD SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_DCAPX1_CV.sym # of pins=2
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DCAPX1_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DCAPX1_CV.sch
.subckt SUNTR_DCAPX1_CV A B
*.iopin A
*.iopin B
R1 A NC0 sky130_fd_pr__res_generic_l1 W=0.44 L=0.36 m=1
R2 B NC1 sky130_fd_pr__res_generic_l1 W=0.44 L=0.36 m=1
.ends


* expanding   symbol:  SUN_TRB_SKY130NM/SUNTRB_NCHDL.sym # of pins=4
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_trb_sky130nm/design/SUN_TRB_SKY130NM/SUNTRB_NCHDL.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_trb_sky130nm/design/SUN_TRB_SKY130NM/SUNTRB_NCHDL.sch
.subckt SUNTRB_NCHDL D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.18 W=1.08 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'  sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  SUN_TRB_SKY130NM/SUNTRB_PCHDL.sym # of pins=4
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_trb_sky130nm/design/SUN_TRB_SKY130NM/SUNTRB_PCHDL.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_trb_sky130nm/design/SUN_TRB_SKY130NM/SUNTRB_PCHDL.sch
.subckt SUNTRB_PCHDL D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.18 W=1.08 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'  pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'  sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NDX1_CV.sym # of pins=5
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NDX1_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NDX1_CV.sch
.subckt SUNTR_NDX1_CV A B Y AVDD AVSS
*.iopin A
*.iopin B
*.iopin Y
*.iopin AVDD
*.iopin AVSS
XMN0 N1 A AVSS AVSS SUNTR_NCHDL
XMN1 Y B N1 AVSS SUNTR_NCHDL
XMP0 Y A AVDD AVDD SUNTR_PCHDL
XMP1 AVDD B Y AVDD SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_IVTRIX1_CV.sym # of pins=6
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVTRIX1_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVTRIX1_CV.sch
.subckt SUNTR_IVTRIX1_CV A C CN Y AVDD AVSS
*.iopin A
*.iopin C
*.iopin CN
*.iopin Y
*.iopin AVDD
*.iopin AVSS
XMN0 N1 A AVSS AVSS SUNTR_NCHDL
XMN1 Y C N1 AVSS SUNTR_NCHDL
XMP0 N2 A AVDD AVDD SUNTR_PCHDL
XMP1 Y CN N2 AVDD SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_NDTRIX1_CV.sym # of pins=7
** sym_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NDTRIX1_CV.sym
** sch_path:
*+ /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NDTRIX1_CV.sch
.subckt SUNTR_NDTRIX1_CV A C CN RN Y AVDD AVSS
*.iopin A
*.iopin C
*.iopin CN
*.iopin RN
*.iopin Y
*.iopin AVDD
*.iopin AVSS
XMN0 N2 A N1 AVSS SUNTR_NCHDL
XMN1 Y C N2 AVSS SUNTR_NCHDL
XMN2 N1 RN AVSS AVSS SUNTR_NCHDL
XMP0 N2 A AVDD AVDD SUNTR_PCHDL
XMP1 Y CN N2 AVDD SUNTR_PCHDL
XMP2 AVDD RN N2 AVDD SUNTR_PCHDL
.ends


* expanding   symbol:  SUN_TR_SKY130NM/SUNTR_RES8.sym # of pins=3
** sym_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RES8.sym
** sch_path: /Users/wulff/data/2023/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RES8.sch
.subckt SUNTR_RES8 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.72 L=8.8 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.72 L=8.8 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.72 L=8.8 mult=1 m=1
XR1_3 INT_3 INT_2 B sky130_fd_pr__res_high_po W=0.72 L=8.8 mult=1 m=1
XR1_4 INT_4 INT_3 B sky130_fd_pr__res_high_po W=0.72 L=8.8 mult=1 m=1
XR1_5 INT_5 INT_4 B sky130_fd_pr__res_high_po W=0.72 L=8.8 mult=1 m=1
XR1_6 INT_6 INT_5 B sky130_fd_pr__res_high_po W=0.72 L=8.8 mult=1 m=1
XR1_7 P INT_6 B sky130_fd_pr__res_high_po W=0.72 L=8.8 mult=1 m=1
.ends

.end
