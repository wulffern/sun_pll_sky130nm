* NGSPICE file created from SUN_PLL_ROSC.ext - technology: sky130B

.subckt SUNTRB_PCHDL D G S B a_216_n18# a_216_334# VSUBS
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
C0 a_216_n18# B 0.331f
C1 a_216_334# B 0.331f
C2 B G 0.339f
C3 B VSUBS 2.81f
.ends

.subckt SUNTRB_NCHDL D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
C0 G B 0.412f
C1 a_324_n18# B 0.422f
C2 a_324_334# B 0.422f
.ends

.subckt SUNTRB_IVX1_CV BULKP AVDD AVSS A Y MP0/a_216_n18# MP0/a_216_334# MN0/a_324_n18#
+ VSUBS MN0/a_324_334#
XMP0 Y A AVDD BULKP MP0/a_216_n18# MP0/a_216_334# VSUBS SUNTRB_PCHDL
XMN0 Y A AVSS VSUBS MN0/a_324_n18# MN0/a_324_334# SUNTRB_NCHDL
C0 BULKP A 0.109f
C1 AVSS VSUBS 0.356f
C2 Y VSUBS 0.264f
C3 MN0/a_324_n18# VSUBS 0.422f
C4 MN0/a_324_334# VSUBS 0.422f
C5 AVDD VSUBS 0.245f
C6 A VSUBS 0.628f
C7 BULKP VSUBS 2.81f
.ends

.subckt SUNTRB_NDX1_CV B Y AVDD AVSS MN1/a_324_334# A BULKP MP1/a_216_334# VSUBS
XMP0 Y A AVDD BULKP MP0/a_216_n18# MP1/a_216_n18# VSUBS SUNTRB_PCHDL
XMP1 AVDD B Y BULKP MP1/a_216_n18# MP1/a_216_334# VSUBS SUNTRB_PCHDL
XMN0 MN1/S A AVSS VSUBS MN0/a_324_n18# MN1/a_324_n18# SUNTRB_NCHDL
XMN1 Y B MN1/S VSUBS MN1/a_324_n18# MN1/a_324_334# SUNTRB_NCHDL
C0 BULKP AVDD 0.175f
C1 BULKP MP1/a_216_n18# -0.311f
C2 BULKP Y 0.115f
C3 BULKP B 0.11f
C4 BULKP A 0.11f
C5 AVSS VSUBS 0.411f
C6 MN1/a_324_334# VSUBS 0.422f
C7 AVDD VSUBS 0.345f
C8 MN0/a_324_n18# VSUBS 0.422f
C9 MN1/a_324_n18# VSUBS 0.352f
C10 Y VSUBS 0.299f
C11 B VSUBS 0.561f
C12 BULKP VSUBS 4.38f
C13 A VSUBS 0.562f
.ends

.subckt SUNTRB_TAPCELLBAVSS_CV MN1/a_324_n18# MP1/B MP1/a_216_n18# AVSS
XMP1 MP1/S MP1/S MP1/S MP1/B MP1/a_216_n18# MP1/a_216_334# AVSS SUNTRB_PCHDL
XMN1 AVSS AVSS AVSS AVSS MN1/a_324_n18# MN1/a_324_334# SUNTRB_NCHDL
C0 AVSS 0 1.07f
C1 MN1/a_324_n18# 0 0.422f
C2 MN1/a_324_334# 0 0.422f
C3 MP1/S 0 0.177f
C4 MP1/B 0 2.81f
.ends

.subckt SUNTR_PCHDL D G S B a_216_n18# a_216_334# VSUBS
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
C0 a_216_n18# B 0.331f
C1 a_216_334# B 0.331f
C2 G B 0.339f
C3 B VSUBS 2.81f
.ends

.subckt SUNTR_NCHDL D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
C0 G B 0.412f
C1 a_324_n18# B 0.422f
C2 a_324_334# B 0.422f
.ends

.subckt SUN_PLL_LSCORE A AVDD AVSS xb2_1/a_324_334# xc2b/a_216_334# YN xc2b/B AN Y
+ VSUBS
Xxc2a xc2b/S Y AVDD xc2b/B xc2a/a_216_n18# xc2b/a_216_n18# VSUBS SUNTR_PCHDL
Xxc2b YN Y xc2b/S xc2b/B xc2b/a_216_n18# xc2b/a_216_334# VSUBS SUNTR_PCHDL
Xxc1a xc1b/S YN AVDD xc2b/B xc1a/a_216_n18# xc1b/a_216_n18# VSUBS SUNTR_PCHDL
Xxc1b Y YN xc1b/S xc2b/B xc1b/a_216_n18# xc2a/a_216_n18# VSUBS SUNTR_PCHDL
Xxb1_0 Y AN AVSS VSUBS xb1_0/a_324_n18# xb1_1/a_324_n18# SUNTR_NCHDL
Xxb1_1 Y AN AVSS VSUBS xb1_1/a_324_n18# xb2_0/a_324_n18# SUNTR_NCHDL
Xxb2_0 YN A AVSS VSUBS xb2_0/a_324_n18# xb2_1/a_324_n18# SUNTR_NCHDL
Xxb2_1 YN A AVSS VSUBS xb2_1/a_324_n18# xb2_1/a_324_334# SUNTR_NCHDL
C0 Y AVDD 0.253f
C1 Y AVSS 0.224f
C2 xc2b/a_216_n18# xc2b/B -0.311f
C3 xc2b/B AVDD 0.222f
C4 YN AVSS 0.161f
C5 xc2b/B Y 0.334f
C6 YN Y 0.347f
C7 AVSS AVDD 0.185f
C8 xc1b/a_216_n18# xc2b/B -0.311f
C9 YN xc2b/B 0.414f
C10 xc2a/a_216_n18# xc2b/B -0.311f
C11 AVDD VSUBS 0.362f
C12 AVSS VSUBS 0.742f
C13 xb2_1/a_324_n18# VSUBS 0.352f
C14 xb2_1/a_324_334# VSUBS 0.422f
C15 A VSUBS 0.874f
C16 xb2_0/a_324_n18# VSUBS 0.353f
C17 xb1_1/a_324_n18# VSUBS 0.352f
C18 AN VSUBS 0.874f
C19 Y VSUBS 0.435f
C20 xb1_0/a_324_n18# VSUBS 0.422f
C21 xc2b/B VSUBS 7.54f
C22 YN VSUBS 0.421f
.ends

.subckt SUNTR_IVX1_CV AVDD AVSS MP0/B A Y MP0/a_216_n18# MP0/a_216_334# MN0/a_324_n18#
+ VSUBS MN0/a_324_334#
XMP0 Y A AVDD MP0/B MP0/a_216_n18# MP0/a_216_334# VSUBS SUNTR_PCHDL
XMN0 Y A AVSS VSUBS MN0/a_324_n18# MN0/a_324_334# SUNTR_NCHDL
C0 MP0/B A 0.109f
C1 AVDD VSUBS 0.245f
C2 AVSS VSUBS 0.356f
C3 A VSUBS 0.628f
C4 Y VSUBS 0.264f
C5 MN0/a_324_n18# VSUBS 0.422f
C6 MN0/a_324_334# VSUBS 0.422f
C7 MP0/B VSUBS 2.81f
.ends

.subckt SUNTR_TAPCELLB_CV AVDD MN1/a_324_n18# MP1/a_216_n18# AVSS
XMP1 AVDD AVDD AVDD AVDD MP1/a_216_n18# MP1/a_216_334# AVSS SUNTR_PCHDL
XMN1 AVSS AVSS AVSS AVSS MN1/a_324_n18# MN1/a_324_334# SUNTR_NCHDL
C0 AVDD AVSS 0.105f
C1 AVSS 0 1.04f
C2 MN1/a_324_n18# 0 0.422f
C3 MN1/a_324_334# 0 0.422f
C4 AVDD 0 3.14f
.ends

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt SUN_PLL_ROSC AVDD CK VDD_ROSC PWRUP_1V8 AVSS
*.subckt SUN_PLL_ROSC AVDD CK VDD_ROSC PWRUP_1V8 AVSS
Xxb2_3 AVDD VDD_ROSC AVSS xb2_3/A xb2_4/A xb2_3/MP0/a_216_n18# xb2_4/MP0/a_216_n18#
+ xb2_3/MN0/a_324_n18# AVSS xb2_4/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_2 AVDD VDD_ROSC AVSS xb2_2/A xb2_3/A xb2_2/MP0/a_216_n18# xb2_3/MP0/a_216_n18#
+ xb2_2/MN0/a_324_n18# AVSS xb2_3/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_4 AVDD VDD_ROSC AVSS xb2_4/A xb2_5/A xb2_4/MP0/a_216_n18# xb2_5/MP0/a_216_n18#
+ xb2_4/MN0/a_324_n18# AVSS xb2_5/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_5 AVDD VDD_ROSC AVSS xb2_5/A xa3/A xb2_5/MP0/a_216_n18# xb2_6/MP0/a_216_n18#
+ xb2_5/MN0/a_324_n18# AVSS xb2_6/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_6 AVDD VDD_ROSC AVSS xa3/A xa3/AN xb2_6/MP0/a_216_n18# xb2_7/MP0/a_216_n18# xb2_6/MN0/a_324_n18#
+ AVSS xb2_7/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_7 AVDD VDD_ROSC AVSS xa3/AN xb1/B xb2_7/MP0/a_216_n18# xb3/MP1/a_216_n18# xb2_7/MN0/a_324_n18#
+ AVSS xb3/MN1/a_324_n18# SUNTRB_IVX1_CV
Xxb1 xb1/B xb1/Y VDD_ROSC AVSS xb1/MN1/a_324_334# PWRUP_1V8 AVDD xb1/MP1/a_216_334#
+ AVSS SUNTRB_NDX1_CV
Xxb3 xb3/MN1/a_324_n18# AVDD xb3/MP1/a_216_n18# AVSS SUNTRB_TAPCELLBAVSS_CV
Xxa3 xa3/A AVDD AVSS xa4/MN0/a_324_n18# xa4/MP0/a_216_n18# xa5/A AVDD xa3/AN xa4/A
+ AVSS SUN_PLL_LSCORE
Xxa4 AVDD AVSS AVDD xa4/A xa4/Y xa4/MP0/a_216_n18# xa5/MP0/a_216_n18# xa4/MN0/a_324_n18#
+ AVSS xa5/MN0/a_324_n18# SUNTR_IVX1_CV
Xxa5 AVDD AVSS AVDD xa5/A CK xa5/MP0/a_216_n18# xa6/MP1/a_216_n18# xa5/MN0/a_324_n18#
+ AVSS xa6/MN1/a_324_n18# SUNTR_IVX1_CV
Xxa6 AVDD xa6/MN1/a_324_n18# xa6/MP1/a_216_n18# AVSS SUNTR_TAPCELLB_CV
Xxb2_0 AVDD VDD_ROSC AVSS xb1/Y xb2_1/A xb1/MP1/a_216_334# xb2_1/MP0/a_216_n18# xb1/MN1/a_324_334#
+ AVSS xb2_1/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_1 AVDD VDD_ROSC AVSS xb2_1/A xb2_2/A xb2_1/MP0/a_216_n18# xb2_2/MP0/a_216_n18#
+ xb2_1/MN0/a_324_n18# AVSS xb2_2/MN0/a_324_n18# SUNTRB_IVX1_CV
C0 xa5/A xa4/A 0.241f
C1 AVDD CK 0.436f
C2 xb2_6/MP0/a_216_n18# AVDD -0.311f
C3 VDD_ROSC xa3/A 0.305f
C4 xb2_7/MP0/a_216_n18# AVDD -0.311f
C5 xa6/MP1/a_216_n18# AVDD -0.311f
C6 xa5/A AVDD 0.115f
C7 xb3/MP1/a_216_n18# AVDD -0.311f
C8 VDD_ROSC xa3/AN 0.302f
C9 xb2_2/A xb2_1/A 0.134f
C10 xb2_4/A xb2_5/A 0.134f
C11 xa3/AN xa3/A 0.957f
C12 xa4/A xa3/A 0.288f
C13 xb1/B xa3/AN 0.131f
C14 xb2_4/MP0/a_216_n18# AVDD -0.31f
C15 xa5/MP0/a_216_n18# AVDD -0.311f
C16 xa4/A xa3/AN 0.121f
C17 xb2_5/MP0/a_216_n18# AVDD -0.31f
C18 xb1/B xb1/Y 0.112f
C19 xa4/MP0/a_216_n18# AVDD -0.311f
C20 xb2_5/A xa3/A 0.165f
C21 VDD_ROSC AVDD 0.154f
C22 AVDD xa3/A 0.406f
C23 xb2_3/MP0/a_216_n18# AVDD -0.31f
C24 xb2_1/A xb1/Y 0.121f
C25 xb2_2/MP0/a_216_n18# AVDD -0.31f
C26 xb2_3/A xb2_4/A 0.134f
C27 AVDD xb2_1/MP0/a_216_n18# -0.31f
C28 AVDD xa3/AN 0.283f
C29 xb1/MP1/a_216_334# AVDD -0.31f
C30 AVDD xa4/A 0.103f
C31 PWRUP_1V8 AVDD 0.302f
C32 xb2_3/A xb2_2/A 0.134f
C33 xb2_1/MN0/a_324_n18# AVSS 0.352f
C34 xb2_1/A AVSS 0.786f
C35 xb1/Y AVSS 0.92f
C36 xa6/MN1/a_324_n18# AVSS 0.354f
C37 xa6/MN1/a_324_334# AVSS 0.422f
C38 CK AVSS 1.57f
C39 xa5/MN0/a_324_n18# AVSS 0.356f
C40 xa4/Y AVSS 0.319f
C41 xa4/MN0/a_324_n18# AVSS 0.352f
C42 xa3/xb2_1/a_324_n18# AVSS 0.355f
C43 xa3/A AVSS 3.01f
C44 xa3/xb2_0/a_324_n18# AVSS 0.355f
C45 xa3/xb1_1/a_324_n18# AVSS 0.352f
C46 xa3/AN AVSS 2.99f
C47 xa4/A AVSS 1.57f
C48 xa3/xb1_0/a_324_n18# AVSS 0.467f
C49 AVDD AVSS 36.8f
C50 xa5/A AVSS 1.15f
C51 xa3/xc1a/a_216_n18# AVSS 0.13f
C52 xb3/MN1/a_324_334# AVSS 0.461f
C53 xb3/MP1/S AVSS 0.233f
C54 xb3/MP1/a_216_334# AVSS 0.129f
C55 xb1/MN1/a_324_334# AVSS 0.353f
C56 VDD_ROSC AVSS 0.785f
C57 xb1/MN0/a_324_n18# AVSS 0.469f
C58 xb1/MN1/a_324_n18# AVSS 0.358f
C59 xb1/B AVSS 2.5f
C60 PWRUP_1V8 AVSS 1.23f
C61 xb1/MP0/a_216_n18# AVSS 0.131f
C62 xb3/MN1/a_324_n18# AVSS 0.354f
C63 xb2_6/MN0/a_324_n18# AVSS 0.349f
C64 xb2_7/MN0/a_324_n18# AVSS 0.349f
C65 xb2_5/MN0/a_324_n18# AVSS 0.352f
C66 xb2_5/A AVSS 0.782f
C67 xb2_4/MN0/a_324_n18# AVSS 0.352f
C68 xb2_4/A AVSS 0.782f
C69 xb2_2/MN0/a_324_n18# AVSS 0.352f
C70 xb2_2/A AVSS 0.782f
C71 xb2_3/MN0/a_324_n18# AVSS 0.352f
C72 xb2_3/A AVSS 0.782f
.ends

