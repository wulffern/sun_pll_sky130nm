magic
tech sky130B
magscale 1 1
timestamp 1720908000
<< checkpaint >>
rect 0 0 5952 6328
<< locali >>
rect 5640 192 5760 6120
rect 192 192 5760 312
rect 192 6000 5760 6120
rect 192 192 312 6120
rect 5640 192 5760 6120
rect 5832 0 5952 6312
rect 0 0 5952 120
rect 0 6192 5952 6312
rect 0 0 120 6312
rect 5832 0 5952 6312
rect 816 1205 900 1235
rect 816 1293 900 1323
rect 816 2173 900 2203
rect 816 3053 900 3083
rect 816 3933 900 3963
rect 900 1205 930 3963
rect 585 3097 615 4007
rect 585 1337 615 2247
rect 1662 457 1746 487
rect 1662 721 1746 751
rect 1662 985 1746 1015
rect 1662 1249 1746 1279
rect 1662 1513 1746 1543
rect 1662 1777 1746 1807
rect 1662 2041 1746 2071
rect 1662 2305 1746 2335
rect 1662 2569 1746 2599
rect 1662 2833 1746 2863
rect 1662 3097 1746 3127
rect 1662 3361 1746 3391
rect 1662 3625 1746 3655
rect 1662 3889 1746 3919
rect 1662 4153 1746 4183
rect 1662 4417 1746 4447
rect 1662 4681 1746 4711
rect 1662 4945 1746 4975
rect 1662 5209 1746 5239
rect 1662 5473 1746 5503
rect 1662 5737 1746 5767
rect 1746 457 1776 5767
<< m1 >>
rect 762 192 870 443
rect 330 192 438 494
rect 1608 0 1716 487
rect 1176 0 1284 538
rect 1446 5781 1530 5811
rect 816 4725 1530 4755
rect 1530 1601 1662 1631
rect 1530 1865 1662 1895
rect 1530 2129 1662 2159
rect 1530 2393 1662 2423
rect 1446 2613 1530 2643
rect 1446 2877 1530 2907
rect 1446 3141 1530 3171
rect 1446 3405 1530 3435
rect 1446 3669 1530 3699
rect 1446 3933 1530 3963
rect 1446 4197 1530 4227
rect 1446 4461 1530 4491
rect 1446 4725 1530 4755
rect 1446 4989 1530 5019
rect 1446 5253 1530 5283
rect 1446 5517 1530 5547
rect 816 3845 1530 3875
rect 1530 1601 1560 5811
rect 0 3097 108 3127
rect 0 3097 108 3127
rect 486 3097 600 3127
rect 54 3097 486 3127
rect 486 3097 516 3127
<< m3 >>
rect 3714 192 3822 404
rect 1662 2657 1752 2695
rect 1662 2921 1752 2959
rect 1662 3185 1752 3223
rect 1662 3449 1752 3487
rect 1662 3713 1752 3751
rect 1662 3977 1752 4015
rect 1662 4241 1752 4279
rect 1662 4505 1752 4543
rect 1662 4769 1752 4807
rect 1662 5033 1752 5071
rect 1662 5297 1752 5335
rect 1662 5561 1752 5599
rect 1662 5825 1752 5863
rect 1752 764 3768 802
rect 1752 1244 3768 1282
rect 1752 1724 3768 1762
rect 1752 2204 3768 2242
rect 1752 2684 3768 2722
rect 1752 3164 3768 3202
rect 1752 3644 3768 3682
rect 1752 4124 3768 4162
rect 1752 4604 3768 4642
rect 1752 5084 3768 5122
rect 1752 5564 3768 5602
rect 1752 764 1790 5863
rect 3768 364 5694 402
rect 3768 844 5694 882
rect 3768 1324 5694 1362
rect 3768 1804 5694 1842
rect 3768 2284 5694 2322
rect 3768 2764 5694 2802
rect 3768 3244 5694 3282
rect 3768 3724 5694 3762
rect 3768 4204 5694 4242
rect 3768 4684 5694 4722
rect 3768 5164 5694 5202
rect 5694 364 5732 5202
rect 546 6282 654 6312
rect 1608 6290 1716 6320
rect 546 6282 654 6312
rect 472 1337 600 1375
rect 472 6282 600 6320
rect 472 1337 510 6320
rect 1608 6290 1716 6320
rect 1662 2657 1752 2695
rect 1662 6290 1752 6328
rect 1752 2657 1790 6328
<< m2 >>
rect 1446 501 1532 539
rect 816 2965 1532 3003
rect 1532 545 1662 583
rect 816 2085 1532 2123
rect 1532 809 1662 847
rect 1446 765 1532 803
rect 1532 1073 1662 1111
rect 1446 1029 1532 1067
rect 1532 1337 1662 1375
rect 1446 1293 1532 1331
rect 1446 1557 1532 1595
rect 1446 1821 1532 1859
rect 1446 2085 1532 2123
rect 1446 2349 1532 2387
rect 1532 501 1570 3003
rect 0 457 108 487
rect 0 457 108 487
rect 476 457 600 495
rect 54 457 476 495
rect 476 457 514 495
use SUNTR_NCHDLCM xa1 ../SUN_TR_SKY130NM
transform 1 0 384 0 1 384
box 384 384 1014 1264
use SUNTR_NCHDLCM xa2_0 ../SUN_TR_SKY130NM
transform 1 0 384 0 1 1264
box 384 1264 1014 2144
use SUNTR_NCHDLCM xa2_1 ../SUN_TR_SKY130NM
transform 1 0 384 0 1 2144
box 384 2144 1014 3024
use SUNTR_NCHDLCM xa4_0 ../SUN_TR_SKY130NM
transform 1 0 384 0 1 3024
box 384 3024 1014 3904
use SUNTR_NCHDLCM xa4_1 ../SUN_TR_SKY130NM
transform 1 0 384 0 1 3904
box 384 3904 1014 4784
use SUNTR_PCHL xc1_0 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 384
box 1860 384 2490 648
use SUNTR_PCHL xc1_1 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 648
box 1860 648 2490 912
use SUNTR_PCHL xc1_2 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 912
box 1860 912 2490 1176
use SUNTR_PCHL xc1_3 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 1176
box 1860 1176 2490 1440
use SUNTR_PCHL xc2_0 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 1440
box 1860 1440 2490 1704
use SUNTR_PCHL xc2_1 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 1704
box 1860 1704 2490 1968
use SUNTR_PCHL xc2_2 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 1968
box 1860 1968 2490 2232
use SUNTR_PCHL xc2_3 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 2232
box 1860 2232 2490 2496
use SUNTR_PCHL xc3_0 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 2496
box 1860 2496 2490 2760
use SUNTR_PCHL xc3_1 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 2760
box 1860 2760 2490 3024
use SUNTR_PCHL xc3_10 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 3024
box 1860 3024 2490 3288
use SUNTR_PCHL xc3_11 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 3288
box 1860 3288 2490 3552
use SUNTR_PCHL xc3_12 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 3552
box 1860 3552 2490 3816
use SUNTR_PCHL xc3_2 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 3816
box 1860 3816 2490 4080
use SUNTR_PCHL xc3_3 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 4080
box 1860 4080 2490 4344
use SUNTR_PCHL xc3_4 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 4344
box 1860 4344 2490 4608
use SUNTR_PCHL xc3_5 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 4608
box 1860 4608 2490 4872
use SUNTR_PCHL xc3_6 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 4872
box 1860 4872 2490 5136
use SUNTR_PCHL xc3_7 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 5136
box 1860 5136 2490 5400
use SUNTR_PCHL xc3_8 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 5400
box 1860 5400 2490 5664
use SUNTR_PCHL xc3_9 ../SUN_TR_SKY130NM
transform -1 0 1860 0 1 5664
box 1860 5664 2490 5928
use SUNSAR_CAP_BSSW_CV xd2 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 384
box 1932 384 5568 864
use SUNSAR_CAP_BSSW_CV xd3_0 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 864
box 1932 864 5568 1344
use SUNSAR_CAP_BSSW_CV xd3_1 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 1344
box 1932 1344 5568 1824
use SUNSAR_CAP_BSSW_CV xd3_2 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 1824
box 1932 1824 5568 2304
use SUNSAR_CAP_BSSW_CV xd3_3 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 2304
box 1932 2304 5568 2784
use SUNSAR_CAP_BSSW_CV xd3_4 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 2784
box 1932 2784 5568 3264
use SUNSAR_CAP_BSSW_CV xd3_5 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 3264
box 1932 3264 5568 3744
use SUNSAR_CAP_BSSW_CV xd3_6 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 3744
box 1932 3744 5568 4224
use SUNSAR_CAP_BSSW_CV xd3_7 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 4224
box 1932 4224 5568 4704
use SUNSAR_CAP_BSSW_CV xd3_8 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 4704
box 1932 4704 5568 5184
use SUNSAR_CAP_BSSW_CV xd3_9 ../SUN_SAR9B_SKY130NM
transform 1 0 1932 0 1 5184
box 1932 5184 5568 5664
use cut_M1M2_2x1 xcut0 
transform 1 0 770 0 1 413
box 770 413 862 447
use cut_M1M2_2x1 xcut1 
transform 1 0 770 0 1 192
box 770 192 862 226
use cut_M1M2_2x1 xcut2 
transform 1 0 338 0 1 450
box 338 450 430 484
use cut_M1M2_2x1 xcut3 
transform 1 0 338 0 1 192
box 338 192 430 226
use cut_M1M4_2x1 xcut4 
transform 1 0 3718 0 1 192
box 3718 192 3818 230
use cut_M1M2_2x1 xcut5 
transform 1 0 1616 0 1 457
box 1616 457 1708 491
use cut_M1M2_2x1 xcut6 
transform 1 0 1616 0 1 0
box 1616 0 1708 34
use cut_M1M2_2x1 xcut7 
transform 1 0 1184 0 1 494
box 1184 494 1276 528
use cut_M1M2_2x1 xcut8 
transform 1 0 1184 0 1 0
box 1184 0 1276 34
use cut_M1M2_2x1 xcut9 
transform 1 0 1392 0 1 5781
box 1392 5781 1484 5815
use cut_M1M2_2x1 xcut10 
transform 1 0 762 0 1 4725
box 762 4725 854 4759
use cut_M1M2_2x1 xcut11 
transform 1 0 1608 0 1 1601
box 1608 1601 1700 1635
use cut_M1M2_2x1 xcut12 
transform 1 0 1608 0 1 1865
box 1608 1865 1700 1899
use cut_M1M2_2x1 xcut13 
transform 1 0 1608 0 1 2129
box 1608 2129 1700 2163
use cut_M1M2_2x1 xcut14 
transform 1 0 1608 0 1 2393
box 1608 2393 1700 2427
use cut_M1M2_2x1 xcut15 
transform 1 0 1392 0 1 2613
box 1392 2613 1484 2647
use cut_M1M2_2x1 xcut16 
transform 1 0 1392 0 1 2877
box 1392 2877 1484 2911
use cut_M1M2_2x1 xcut17 
transform 1 0 1392 0 1 3141
box 1392 3141 1484 3175
use cut_M1M2_2x1 xcut18 
transform 1 0 1392 0 1 3405
box 1392 3405 1484 3439
use cut_M1M2_2x1 xcut19 
transform 1 0 1392 0 1 3669
box 1392 3669 1484 3703
use cut_M1M2_2x1 xcut20 
transform 1 0 1392 0 1 3933
box 1392 3933 1484 3967
use cut_M1M2_2x1 xcut21 
transform 1 0 1392 0 1 4197
box 1392 4197 1484 4231
use cut_M1M2_2x1 xcut22 
transform 1 0 1392 0 1 4461
box 1392 4461 1484 4495
use cut_M1M2_2x1 xcut23 
transform 1 0 1392 0 1 4725
box 1392 4725 1484 4759
use cut_M1M2_2x1 xcut24 
transform 1 0 1392 0 1 4989
box 1392 4989 1484 5023
use cut_M1M2_2x1 xcut25 
transform 1 0 1392 0 1 5253
box 1392 5253 1484 5287
use cut_M1M2_2x1 xcut26 
transform 1 0 1392 0 1 5517
box 1392 5517 1484 5551
use cut_M1M2_2x1 xcut27 
transform 1 0 762 0 1 3845
box 762 3845 854 3879
use cut_M1M3_2x1 xcut28 
transform 1 0 1392 0 1 501
box 1392 501 1492 539
use cut_M1M3_2x1 xcut29 
transform 1 0 762 0 1 2965
box 762 2965 862 3003
use cut_M1M3_2x1 xcut30 
transform 1 0 1608 0 1 545
box 1608 545 1708 583
use cut_M1M3_2x1 xcut31 
transform 1 0 762 0 1 2085
box 762 2085 862 2123
use cut_M1M3_2x1 xcut32 
transform 1 0 1608 0 1 809
box 1608 809 1708 847
use cut_M1M3_2x1 xcut33 
transform 1 0 1392 0 1 765
box 1392 765 1492 803
use cut_M1M3_2x1 xcut34 
transform 1 0 1608 0 1 1073
box 1608 1073 1708 1111
use cut_M1M3_2x1 xcut35 
transform 1 0 1392 0 1 1029
box 1392 1029 1492 1067
use cut_M1M3_2x1 xcut36 
transform 1 0 1608 0 1 1337
box 1608 1337 1708 1375
use cut_M1M3_2x1 xcut37 
transform 1 0 1392 0 1 1293
box 1392 1293 1492 1331
use cut_M1M3_2x1 xcut38 
transform 1 0 1392 0 1 1557
box 1392 1557 1492 1595
use cut_M1M3_2x1 xcut39 
transform 1 0 1392 0 1 1821
box 1392 1821 1492 1859
use cut_M1M3_2x1 xcut40 
transform 1 0 1392 0 1 2085
box 1392 2085 1492 2123
use cut_M1M3_2x1 xcut41 
transform 1 0 1392 0 1 2349
box 1392 2349 1492 2387
use cut_M1M4_2x1 xcut42 
transform 1 0 1608 0 1 2657
box 1608 2657 1708 2695
use cut_M1M4_2x1 xcut43 
transform 1 0 1608 0 1 2921
box 1608 2921 1708 2959
use cut_M1M4_2x1 xcut44 
transform 1 0 1608 0 1 3185
box 1608 3185 1708 3223
use cut_M1M4_2x1 xcut45 
transform 1 0 1608 0 1 3449
box 1608 3449 1708 3487
use cut_M1M4_2x1 xcut46 
transform 1 0 1608 0 1 3713
box 1608 3713 1708 3751
use cut_M1M4_2x1 xcut47 
transform 1 0 1608 0 1 3977
box 1608 3977 1708 4015
use cut_M1M4_2x1 xcut48 
transform 1 0 1608 0 1 4241
box 1608 4241 1708 4279
use cut_M1M4_2x1 xcut49 
transform 1 0 1608 0 1 4505
box 1608 4505 1708 4543
use cut_M1M4_2x1 xcut50 
transform 1 0 1608 0 1 4769
box 1608 4769 1708 4807
use cut_M1M4_2x1 xcut51 
transform 1 0 1608 0 1 5033
box 1608 5033 1708 5071
use cut_M1M4_2x1 xcut52 
transform 1 0 1608 0 1 5297
box 1608 5297 1708 5335
use cut_M1M4_2x1 xcut53 
transform 1 0 1608 0 1 5561
box 1608 5561 1708 5599
use cut_M1M4_2x1 xcut54 
transform 1 0 1608 0 1 5825
box 1608 5825 1708 5863
use cut_M1M3_2x1 xcut55 
transform 1 0 554 0 1 457
box 554 457 654 495
use cut_M1M4_2x1 xcut56 
transform 1 0 554 0 1 1337
box 554 1337 654 1375
use cut_M1M2_2x1 xcut57 
transform 1 0 562 0 1 3097
box 562 3097 654 3131
<< labels >>
flabel locali s 5640 192 5760 6120 0 FreeSans 400 0 0 0 AVSS
port 6 nsew signal bidirectional
flabel locali s 5832 0 5952 6312 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel m3 s 546 6282 654 6312 0 FreeSans 400 0 0 0 VFB
port 2 nsew signal bidirectional
flabel m1 s 0 3097 108 3127 0 FreeSans 400 0 0 0 VI
port 3 nsew signal bidirectional
flabel m3 s 1608 6290 1716 6320 0 FreeSans 400 0 0 0 VO
port 4 nsew signal bidirectional
flabel m2 s 0 457 108 487 0 FreeSans 400 0 0 0 VBN
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 5952 6328
<< end >>
