

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
*.include ../../../work/lpe/SUN_PLL_lpe.spi
.include ../../../work/lpe/SUN_PLL_LPF_lpe.spi
.include ../../../work/lpe/SUN_PLL_BUF_lpe.spi
.include ../../../work/lpe/SUN_PLL_ROSC_lpe.spi
.include ../../../work/lpe/SUN_PLL_DIVN_lpe.spi
.include ../../../work/lpe/SUN_PLL_KICK_lpe.spi
.include ../../../work/lpe/SUN_PLL_PFD_lpe.spi
.include ../../../work/lpe/SUN_PLL_CP_lpe.spi
.include ../../../work/lpe/SUN_PLL_BIAS_lpe.spi
.include ../../../design/SUN_PLL_SKY130NM.spice
#else
.include ../../../design/SUN_PLL_SKY130NM.spice
#else
.include ../../../design/SUN_PLL_SKY130NM.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
#ifdef Debug
.option reltol=1e-3 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-12
#else
.option reltol=1e-5 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-15
#endif

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param PERIOD_CLK = 62.5n
.param PW_CLK = PERIOD_CLK/2

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  AVSS  0     dc 0
VDD  AVDD  AVSS  dc  {AVDD}
VPWR  PWRUP_1V8  AVSS pwl 0 0 10n 0 11n {AVDD}

IDC 0 IBPSR_1U  dc 1u


VCKREF CK_REF 0 dc 0 pulse (0 {AVDD} 0 {TRF} {TRF} {PW_CLK} {PERIOD_CLK})
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT AVDD AVSS PWRUP_1V8 CK_REF CK IBPSR_1U SUN_PLL


*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.probe v(AVDD) v(AVSS) v(PWRUP_1V8) v(CK_REF) v(CK) v(IBPSR_1U)
+ v(XDUT.VDD_ROSC) v(XDUT.CP_UP_N) v(XDUT.CP_DOWN) v(XDUT.VLPF) v(XDUT.CK_FB) v(XDUT.KICK) v(XDUT.VLPFZ)
+ v(XDUT.x1.N*)
#else
.probe v(CK_REF) v(CK) v(XDUT.CK_FB) v(XDUT.VDD_ROSC) v(XDUT.CP_UP_N) v(XDUT.CP_DOWN)  v(IBPSR_1U) v(XDUT.VLPF)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=16
set color0=white
set color1=black
unset askquit

#ifdef Debug
tran 10p 500n 1p
write
quit
#else
tran 10p 8u 1p
write
quit
#endif

.endc

.end


