magic
tech sky130B
timestamp 1681076574
<< locali >>
rect 0 5136 2064 5256
rect 0 120 120 5136
rect 192 4944 1872 5064
rect 192 312 312 4944
rect 762 4813 870 4843
rect 600 4593 732 4623
rect 702 4345 732 4593
rect 762 4549 870 4579
rect 702 4315 792 4345
rect 762 4285 816 4315
rect 762 677 870 707
rect 546 633 654 663
rect 1752 312 1872 4944
rect 192 192 1872 312
rect 1944 120 2064 5136
rect 0 0 2064 120
<< metal1 >>
rect 600 4769 714 4799
rect 684 4579 714 4769
rect 684 4549 816 4579
rect 486 4417 600 4447
rect 486 839 516 4417
rect 600 4241 732 4271
rect 702 4169 732 4241
rect 702 4139 792 4169
rect 762 4109 816 4139
rect 600 4065 732 4095
rect 702 3296 732 4065
rect 702 3266 1302 3296
rect 702 3201 732 3266
rect 702 3171 792 3201
rect 762 3141 816 3171
rect 600 3097 732 3127
rect 702 3025 732 3097
rect 702 2995 792 3025
rect 762 2965 816 2995
rect 600 2921 732 2951
rect 702 2152 732 2921
rect 702 2122 1302 2152
rect 702 2057 732 2122
rect 702 2027 792 2057
rect 762 1997 816 2027
rect 600 1953 732 1983
rect 702 1881 732 1953
rect 702 1851 792 1881
rect 762 1821 816 1851
rect 600 1777 732 1807
rect 702 1008 732 1777
rect 702 978 1302 1008
rect 702 913 732 978
rect 702 883 792 913
rect 762 853 816 883
rect 486 809 600 839
rect 486 707 516 809
rect 486 677 816 707
<< metal3 >>
rect 758 192 866 4872
rect 1154 384 1262 5256
use SUNTR_TAPCELLB_CV  xa1a ../SUN_TR_SKY130NM
timestamp 1681076574
transform 1 0 384 0 1 384
box -90 -66 1350 242
use SUNTR_IVX1_CV  xa1b ../SUN_TR_SKY130NM
timestamp 1681076574
transform 1 0 384 0 1 560
box -90 -66 1350 242
use SUNTR_DCAPX1_CV  xa1capd ../SUN_TR_SKY130NM
timestamp 1680904800
transform 1 0 384 0 1 912
box -54 -22 1314 814
use SUNTR_IVX1_CV  xa1c
timestamp 1681076574
transform 1 0 384 0 1 736
box -90 -66 1350 242
use SUNTR_IVX1_CV  xa2
timestamp 1681076574
transform 1 0 384 0 1 1704
box -90 -66 1350 242
use SUNTR_IVX1_CV  xa3a
timestamp 1681076574
transform 1 0 384 0 1 1880
box -90 -66 1350 242
use SUNTR_DCAPX1_CV  xa3capb
timestamp 1680904800
transform 1 0 384 0 1 2056
box -54 -22 1314 814
use SUNTR_IVX1_CV  xa4
timestamp 1681076574
transform 1 0 384 0 1 2848
box -90 -66 1350 242
use SUNTR_IVX1_CV  xa5a
timestamp 1681076574
transform 1 0 384 0 1 3024
box -90 -66 1350 242
use SUNTR_DCAPX1_CV  xa5capb
timestamp 1680904800
transform 1 0 384 0 1 3200
box -54 -22 1314 814
use SUNTR_IVX1_CV  xa6
timestamp 1681076574
transform 1 0 384 0 1 3992
box -90 -66 1350 242
use SUNTR_IVX1_CV  xa7
timestamp 1681076574
transform 1 0 384 0 1 4168
box -90 -66 1350 242
use SUNTR_NRX1_CV  xa8 ../SUN_TR_SKY130NM
timestamp 1681076574
transform 1 0 384 0 1 4344
box -90 -66 1350 418
use SUNTR_IVX1_CV  xa9
timestamp 1681076574
transform 1 0 384 0 1 4696
box -90 -66 1350 242
use cut_M1M2_2x1  xcut0
timestamp 1680991200
transform 1 0 778 0 1 853
box 0 0 92 34
use cut_M1M2_2x1  xcut1
timestamp 1680991200
transform 1 0 1282 0 1 978
box 0 0 92 34
use cut_M1M2_2x1  xcut2
timestamp 1680991200
transform 1 0 562 0 1 1777
box 0 0 92 34
use cut_M1M2_2x1  xcut3
timestamp 1680991200
transform 1 0 778 0 1 1821
box 0 0 92 34
use cut_M1M2_2x1  xcut4
timestamp 1680991200
transform 1 0 562 0 1 1953
box 0 0 92 34
use cut_M1M2_2x1  xcut5
timestamp 1680991200
transform 1 0 778 0 1 1997
box 0 0 92 34
use cut_M1M2_2x1  xcut6
timestamp 1680991200
transform 1 0 1282 0 1 2122
box 0 0 92 34
use cut_M1M2_2x1  xcut7
timestamp 1680991200
transform 1 0 562 0 1 2921
box 0 0 92 34
use cut_M1M2_2x1  xcut8
timestamp 1680991200
transform 1 0 778 0 1 2965
box 0 0 92 34
use cut_M1M2_2x1  xcut9
timestamp 1680991200
transform 1 0 562 0 1 3097
box 0 0 92 34
use cut_M1M2_2x1  xcut10
timestamp 1680991200
transform 1 0 778 0 1 3141
box 0 0 92 34
use cut_M1M2_2x1  xcut11
timestamp 1680991200
transform 1 0 1282 0 1 3266
box 0 0 92 34
use cut_M1M2_2x1  xcut12
timestamp 1680991200
transform 1 0 562 0 1 4065
box 0 0 92 34
use cut_M1M2_2x1  xcut13
timestamp 1680991200
transform 1 0 778 0 1 4109
box 0 0 92 34
use cut_M1M2_2x1  xcut14
timestamp 1680991200
transform 1 0 562 0 1 4241
box 0 0 92 34
use cut_M1M2_2x1  xcut15
timestamp 1680991200
transform 1 0 546 0 1 4769
box 0 0 92 34
use cut_M1M2_2x1  xcut16
timestamp 1680991200
transform 1 0 762 0 1 4549
box 0 0 92 34
use cut_M1M2_2x1  xcut17
timestamp 1680991200
transform 1 0 546 0 1 809
box 0 0 92 34
use cut_M1M2_2x1  xcut18
timestamp 1680991200
transform 1 0 762 0 1 677
box 0 0 92 34
use cut_M1M2_2x1  xcut19
timestamp 1680991200
transform 1 0 546 0 1 4417
box 0 0 92 34
use cut_M1M4_2x1  xcut20
timestamp 1680991200
transform 1 0 762 0 1 192
box 0 0 100 38
use cut_M1M4_2x1  xcut21
timestamp 1680991200
transform 1 0 762 0 1 1594
box 0 0 100 38
use cut_M1M4_2x1  xcut22
timestamp 1680991200
transform 1 0 762 0 1 2738
box 0 0 100 38
use cut_M1M4_2x1  xcut23
timestamp 1680991200
transform 1 0 762 0 1 3882
box 0 0 100 38
use cut_M1M4_2x1  xcut24
timestamp 1680991200
transform 1 0 1158 0 1 5136
box 0 0 100 38
<< labels >>
flabel locali s 1752 192 1872 5064 0 FreeSans 200 0 0 0 AVSS
port 5 nsew signal bidirectional
flabel locali s 1944 0 2064 5256 0 FreeSans 200 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel locali s 762 4549 870 4579 0 FreeSans 200 0 0 0 KICK
port 2 nsew signal bidirectional
flabel locali s 762 4813 870 4843 0 FreeSans 200 0 0 0 KICK_N
port 3 nsew signal bidirectional
flabel locali s 546 633 654 663 0 FreeSans 200 0 0 0 PWRUP_1V8
port 4 nsew signal bidirectional
flabel locali s 762 677 870 707 0 FreeSans 200 0 0 0 PWRUP_1V8_N
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2064 5256
<< end >>
