magic
tech sky130B
magscale 1 2
timestamp 1680904800
<< checkpaint >>
rect 0 0 200 76
<< m2 >>
rect 0 0 200 76
<< m3 >>
rect 0 0 200 76
<< v2 >>
rect 12 6 188 70
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 200 76
<< end >>
