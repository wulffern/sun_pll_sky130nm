* NGSPICE file created from SUN_PLL.ext - technology: sky130B

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt SUN_PLL AVDD AVSS PWRUP_1V8 CK_REF CK IBPSR_1U
*.subckt SUN_PLL PWRUP_1V8 CK_REF CK IBPSR_1U AVSS AVDD
X0 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R0 xaa4.xa2.M0.G m3_22692_52900# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X1 xaa4.xa1.M6.D IBPSR_1U xaa4.xa1.M5.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X2 xaa1.xa2.M8.D IBPSR_1U xaa1.xa2.M7.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X3 xaa6.xf.XA6.MN0.G xaa6.xf.XA5.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X4 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=63.4 pd=346 as=0.616 ps=3.3 w=1.08 l=0.18
X5 xaa6.xf.XA7.MN1.G PWRUP_1V8 xaa6.xf.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X6 xaa0.xa3.MP0.D xaa0.xa1.MN2.S AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X7 AVDD PWRUP_1V8 xaa6.xd.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X8 xaa6.xe.XA7.MP1.G xaa6.xe.XA7.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X9 xaa6.xd.XA5.MN0.G xaa6.xd.XA7.MP1.G xaa6.xd.XA3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X10 xaa6.xf.XA5.MN0.G xaa6.xf.XA7.MP1.G xaa6.xf.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X11 xaa5.xb2_1.MN0.D xaa5.xb2_0.MN0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X12 xaa4.xa1.M8.D IBPSR_1U xaa4.xa1.M7.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R1 AVSS m3_37748_78364# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X13 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MN1.G xaa6.xe.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X14 xaa5.xb3.MP1.D xaa5.xb3.MP1.D xaa5.xb3.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=1.23 pd=6.6 as=0.616 ps=3.3 w=1.08 l=0.18
R2 m3_4628_81084# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X15 xaa6.xe.XA3.MP0.D xaa6.xe.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X16 xaa6.xd.XA4.MP0.D xaa6.xd.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X17 xaa5.xb2_2.MN0.D xaa5.xb2_1.MN0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X18 a_2084_70022# xaa1.xa3.D AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R3 m3_13116_61524# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X19 xaa6.xe.XA6.MP0.D xaa6.xe.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R4 AVSS m3_37748_73564# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X20 xaa6.xc.XA7.MP1.G xaa6.xc.XA7.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X21 xaa5.xb1.MN1.G xaa5.xa3.xb1_0.G xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X22 xaa1.xa2.M7.D IBPSR_1U xaa1.xa2.M6.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R5 m3_4628_89724# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X23 xaa1.xb2.M0.D xaa1.xa1.M8.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X24 xaa1.xa1.M5.D IBPSR_1U xaa1.xa1.M4.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R6 xaa4.xa2.M0.G m3_22692_61348# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R7 m3_13116_55188# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X25 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MP1.G xaa6.xc.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X26 a_356_74698# a_n76_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X27 xaa1.xa2.M5.D IBPSR_1U xaa1.xa2.M4.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R8 m3_13116_58356# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X28 xaa6.xc.XA3.MN0.D xaa6.xc.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X29 xaa1.xa1.M3.D IBPSR_1U xaa1.xa1.M2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X30 xaa5.xa3.xb2_0.D xaa5.xa3.xb2_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R9 AVSS li_6204_57236# sky130_fd_pr__res_generic_l1 w=0.44 l=0.36
X31 xaa3.xa6.MN0.D xaa3.xa1c.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X32 a_n508_70022# xbb0.xa1.XA1.N AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X33 xaa6.xc.XA6.MN0.D xaa6.xc.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X34 a_2084_74698# a_1652_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R10 m3_4628_84924# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X35 xaa6.xf.XA7.MP1.G xaa6.xf.XA7.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X36 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=59.1 pd=317 as=0.616 ps=3.3 w=1.08 l=0.18
X37 xaa4.xa1.M5.D IBPSR_1U xaa4.xa1.M4.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R11 m3_4628_76284# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X38 xaa6.xd.XA7.MN2.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X39 xaa6.xd.XA5.MN0.G xaa6.xd.XA7.MN1.G xaa6.xd.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X40 xaa5.xb2_1.MN0.D xaa5.xb2_0.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X41 xaa3.xa7.MN0.D xaa3.xa6.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X42 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MN1.G xaa6.xf.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R12 AVSS m3_37748_86044# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X43 xaa4.xa1.M3.D IBPSR_1U xaa4.xa1.M2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X44 xaa6.xf.XA3.MP0.D xaa6.xf.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X45 IBPSR_1U IBPSR_1U xbb1.xa3.M7.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X46 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R13 AVSS m3_37748_89884# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R14 m3_4628_71484# xaa1.xa3.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X47 xaa6.xf.XA6.MP0.D xaa6.xf.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X48 xaa6.xd.XA4.MN0.D xaa6.xd.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X49 xaa5.xa3.xc1a.D xaa5.xa3.xb2_0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X50 xaa5.xb2_2.MN0.D xaa5.xb2_1.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X51 xaa6.xg.XA1.MN0.D CK AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X52 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X53 xaa0.xa1.MN0.D xaa0.xa1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X54 CK xaa5.xa3.xb2_0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X55 xbb1.xa3.M6.D IBPSR_1U xbb1.xa3.M5.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X56 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R15 AVSS m3_37748_81244# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X57 AVDD PWRUP_1V8 xaa6.xg.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X58 xaa5.xb1.MN1.G xaa5.xa3.xb1_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X59 xaa6.xc.XA7.MN1.G xaa6.xc.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X60 xaa6.xe.XA6.MN0.G xaa6.xe.XA5.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X61 xaa6.xg.XA5.MN0.G xaa6.xg.XA7.MP1.G xaa6.xg.XA3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X62 xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X63 xaa6.xe.XA7.MN1.G PWRUP_1V8 xaa6.xe.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X64 xaa4.xa4.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X65 xaa1.xa4.M0.D xaa1.xa4.M0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X66 xaa3.xa1b.MN0.D PWRUP_1V8 AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X67 xaa1.xa2.M0.D IBPSR_1U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X68 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X69 xaa6.xe.XA5.MN0.G xaa6.xe.XA7.MP1.G xaa6.xe.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X70 a_1220_70022# a_1652_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X71 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MN1.G xaa6.xg.XA7.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X72 xaa6.xg.XA4.MP0.D xaa6.xg.XA4.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R16 m3_4628_92604# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X73 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MP1.G xaa6.xc.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X74 xaa6.xf.XA7.MP1.G xaa6.xf.XA7.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X75 xaa4.xa1.M0.D IBPSR_1U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X76 xaa6.xg.XA7.MN0.D xaa6.xg.XA7.MN0.G xaa6.xg.XA7.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X77 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X78 xaa1.xa2.M2.D IBPSR_1U xaa1.xa2.M1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X79 xaa0.xa1.MP1.D xaa0.xa1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R17 xaa4.xa2.M0.G m3_22692_60292# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X80 xaa6.xc.XA7.MN0.D xaa0.xa5.MN2.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R18 xaa4.xa2.M0.G m3_22692_63460# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X81 xaa4.xa2.M0.D xaa4.xa2.M0.G xaa4.xa1.M8.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X82 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MP1.G xaa6.xf.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X83 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R19 AVSS m3_37748_76444# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X84 xaa6.xf.XA3.MN0.D xaa6.xf.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X85 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X86 xaa5.xb1.MN1.D PWRUP_1V8 xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X87 AVDD PWRUP_1V8 xaa6.xe.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X88 xbb1.xa3.M3.D IBPSR_1U xbb1.xa3.M2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X89 xaa6.xe.XA5.MN0.G xaa6.xe.XA7.MP1.G xaa6.xe.XA3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X90 xaa6.xf.XA6.MN0.D xaa6.xf.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X91 xaa5.xb2_3.MN0.D xaa5.xb2_2.MN0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X92 xaa6.xd.XA7.MN1.G xaa6.xd.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X93 xbb1.xa3.M1.D IBPSR_1U xbb1.xa3.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R20 AVSS m3_37748_71644# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R21 m3_13116_54132# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R22 m3_13116_57300# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X94 xaa6.xe.XA4.MP0.D xaa6.xe.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X95 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
R23 m3_4628_87804# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X96 xaa5.xb2_4.MN0.D xaa5.xb2_3.MN0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R24 AVSS m3_37748_92764# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X97 xaa6.xc.XA7.MN2.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R25 m3_4628_79164# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X98 xaa6.xc.XA5.MN0.G xaa6.xc.XA7.MN1.G xaa6.xc.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X99 xaa5.xa3.xb2_0.D xaa5.xa3.xb2_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X100 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MP1.G xaa6.xd.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X101 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
R26 xaa4.xa2.M0.G m3_22692_57124# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X102 xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X103 xaa4.xa4.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X104 xaa6.xd.XA7.MN0.D xaa6.xc.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X105 xaa6.xc.XA4.MN0.D xaa6.xc.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X106 xaa1.xa1.M7.D IBPSR_1U xaa1.xa1.M6.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X107 xaa5.xa4.MN0.D xaa5.xa3.xb1_0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R27 m3_4628_74364# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X108 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X109 AVDD PWRUP_1V8 xaa6.xf.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R28 AVSS m3_37748_84124# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X110 xaa6.xf.XA5.MN0.G xaa6.xf.XA7.MP1.G xaa6.xf.XA3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X111 xaa5.xb1.MN0.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X112 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X113 xaa3.xa8.MP0.D xaa3.xa1b.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X114 IBPSR_1U xaa3.xa1b.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R29 AVSS m3_37748_87964# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X115 xaa5.xb2_3.MN0.D xaa5.xb2_2.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X116 a_356_70022# a_n76_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X117 xaa6.xd.XA1.MN0.D xaa6.xd.XA1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X118 xaa4.xa1.M7.D IBPSR_1U xaa4.xa1.M6.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X119 xaa6.xf.XA4.MP0.D xaa6.xf.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X120 a_356_74698# a_788_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R30 m3_4628_90684# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X121 xaa1.xa4.M0.G xaa3.xa7.MN0.D xaa3.xa8.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X122 a_2084_70022# a_1652_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X123 xaa6.xe.XA7.MP1.G xaa6.xe.XA7.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X124 xaa5.xb2_4.MN0.D xaa5.xb2_3.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X125 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
R31 m3_4628_69564# xaa1.xa3.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X126 xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X127 xaa5.xa3.xb1_0.D xaa5.xa3.xb2_0.D xaa5.xa3.xc1a.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X128 xaa4.xa4.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X129 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MP1.G xaa6.xe.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X130 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MN1.G xaa6.xd.XA7.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X131 xaa6.xf.XA1.MN0.G xaa6.xg.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X132 xaa6.xg.XA3.MN1.G CK AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X133 xaa6.xe.XA3.MN0.D xaa6.xe.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X134 xaa6.xg.XA5.MN0.D xaa6.xg.XA5.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R32 AVSS m3_37748_79324# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X135 xaa0.xa5.MN0.D xaa0.xa1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X136 xaa0.xa5.MN2.G xaa6.xc.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X137 xaa6.xg.XA3.MN1.G PWRUP_1V8 xaa6.xg.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X138 a_n508_74698# a_n76_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X139 xaa6.xc.XA6.MN0.G xaa6.xc.XA5.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R33 m3_13116_60468# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X140 xaa0.xa1.MN2.D CK_REF xaa0.xa1.MN2.S AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X141 xaa6.xe.XA6.MN0.D xaa6.xe.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X142 xaa6.xd.XA7.MN0.D xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R34 m3_13116_63636# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X143 AVDD PWRUP_1V8 xaa6.xc.XA7.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R35 m3_4628_82044# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X144 xaa6.xg.XA5.MN0.G xaa6.xg.XA7.MP1.G xaa6.xg.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X145 xaa1.xa1.M2.D IBPSR_1U xaa1.xa1.M1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X146 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X147 AVSS xaa0.xa3.MN1.G xaa0.xa1.MN0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X148 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X149 xaa6.xf.XA7.MN2.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X150 xaa6.xc.XA5.MN0.G xaa6.xc.XA7.MN1.G xaa6.xc.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R36 m3_4628_85884# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X151 xaa6.xf.XA5.MN0.G xaa6.xf.XA7.MN1.G xaa6.xf.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X152 xaa3.xa1b.MN0.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R37 AVSS m3_37748_74524# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X153 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MP1.G xaa6.xg.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X154 xbb1.xa3.M5.D IBPSR_1U xbb1.xa3.M4.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X155 xaa4.xa1.M2.D IBPSR_1U xaa4.xa1.M1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X156 xaa6.xg.XA7.MN0.D xaa6.xg.XA7.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X157 xaa6.xf.XA4.MN0.D xaa6.xf.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X158 xaa0.xa5.MP1.D xaa0.xa1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X159 xbb1.xa3.M7.D IBPSR_1U xbb1.xa3.M6.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X160 xaa0.xa1.MN0.D CK_REF xaa0.xa1.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X161 xaa6.xe.XA7.MN1.G xaa6.xe.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X162 xaa3.xa1c.MN0.D xaa3.xa1b.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X163 xaa4.xa2.M0.G xaa5.xb1.MN1.G xaa5.xb1.MN1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X164 xaa0.xa1.MN0.G xaa0.xa3.MN1.G xaa0.xa3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R38 AVSS m3_37748_90844# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R39 m3_4628_77244# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X165 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X166 xaa6.xd.XA6.MN0.G xaa6.xd.XA5.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X167 xaa5.xa3.xb1_0.D xaa5.xa3.xb1_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R40 AVSS m3_37748_87004# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X168 AVDD PWRUP_1V8 xaa6.xd.XA7.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R41 AVSS m3_37748_69724# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X169 CK xaa5.xa3.xb2_0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X170 xaa4.xa2.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X171 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MP1.G xaa6.xe.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X172 xaa6.xd.XA5.MN0.G xaa6.xd.XA7.MN1.G xaa6.xd.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X173 xaa6.xc.XA1.MN0.D xaa6.xc.XA1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R42 m3_4628_72444# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X174 xaa6.xe.XA7.MN0.D xaa6.xd.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R43 AVSS m3_37748_82204# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X175 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X176 a_1220_74698# a_788_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R44 m3_13116_62580# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X177 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MN1.G xaa6.xc.XA7.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X178 xaa6.xf.XA7.MN1.G xaa6.xf.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X179 xaa3.xa9.MN0.D xaa1.xa4.M0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X180 xbb1.xa3.M2.D IBPSR_1U xbb1.xa3.M1.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X181 xaa1.xb1.M0.D xaa1.xa1.M8.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X182 xaa6.xc.XA7.MN0.D xaa0.xa5.MN2.G xaa6.xc.XA7.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X183 xaa5.xb1.MN1.D xaa5.xb1.MN1.G xaa5.xb1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X184 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X185 xbb1.xa3.M0.D IBPSR_1U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X186 xaa6.xe.XA7.MN2.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X187 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X188 xaa1.xa4.M0.G xaa3.xa1b.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X189 xaa1.xa1.M0.D IBPSR_1U AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X190 xaa6.xe.XA5.MN0.G xaa6.xe.XA7.MN1.G xaa6.xe.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X191 xaa6.xd.XA6.MN0.G xaa6.xd.XA5.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R45 m3_4628_88764# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X192 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MP1.G xaa6.xf.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X193 xaa6.xd.XA7.MN1.G PWRUP_1V8 xaa6.xd.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X194 xaa6.xg.XA7.MP1.G xaa6.xg.XA3.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R46 AVSS m3_37748_77404# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X195 AVSS xaa0.xa1.MN0.D xaa0.xa1.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X196 xaa6.xc.XA7.MP1.G xaa6.xc.XA7.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X197 xaa6.xd.XA5.MN0.G xaa6.xd.XA7.MP1.G xaa6.xd.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X198 AVSS xaa3.xa7.MN0.D xaa1.xa4.M0.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R47 m3_4628_80124# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X199 xaa6.xf.XA7.MN0.D xaa6.xe.XA1.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X200 xaa6.xe.XA4.MN0.D xaa6.xe.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X201 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MP1.G xaa6.xg.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R48 m3_13116_53076# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R49 xaa4.xa2.M0.G m3_22692_62404# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X202 AVSS xaa0.xa5.MN0.D xaa0.xa5.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X203 a_356_70022# a_788_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R50 m3_13116_56244# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X204 xaa6.xg.XA3.MN0.D xaa6.xg.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R51 m3_13116_59412# AVSS sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R52 m3_4628_83964# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X205 xaa0.xa2a.MN0.G xaa0.xa1.MN2.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X206 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MN1.G xaa6.xc.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X207 xaa6.xf.XA1.MN0.G xaa6.xg.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R53 AVSS m3_37748_72604# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X208 xaa6.xc.XA3.MP0.D xaa6.xc.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X209 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X210 xaa6.xg.XA6.MN0.D xaa6.xg.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X211 xaa5.xa3.xc2a.D xaa5.xa3.xb1_0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X212 xaa6.xg.XA5.MN0.D xaa6.xg.XA5.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X213 xaa0.xa5.MN2.D xaa0.xa5.MN2.G xaa0.xa3.MN1.G AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X214 xaa1.xb2.M7.D xaa1.xa1.M8.D xaa1.xb2.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X215 AVDD PWRUP_1V8 xaa6.xg.XA3.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X216 xaa6.xc.XA6.MP0.D xaa6.xc.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R54 xaa4.xa2.M0.G m3_22692_56068# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R55 AVSS m3_37748_85084# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R56 xaa4.xa2.M0.G m3_22692_59236# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X217 xaa1.xa2.M6.D IBPSR_1U xaa1.xa2.M5.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X218 xaa6.xg.XA5.MN0.G xaa6.xg.XA4.MP1.G xaa6.xg.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X219 xaa6.xf.XA1.MN0.D xaa6.xf.XA1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X220 xaa0.xa1.MN2.S xaa0.xa1.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X221 xaa1.xa1.M4.D IBPSR_1U xaa1.xa1.M3.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X222 a_n508_70022# a_n76_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X223 xaa1.xa2.M4.D IBPSR_1U xaa1.xa2.M3.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X224 xaa0.xa3.MN1.G xaa0.xa5.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X225 a_2084_74698# xaa1.xa4.M0.D AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
R57 m3_4628_75324# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X226 xaa4.xa4.M0.D xaa4.xa2.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X227 xaa0.xa2a.MN0.G xaa0.xa1.MN2.S AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R58 AVSS m3_37748_80284# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X228 xaa6.xd.XA7.MP1.G xaa6.xd.XA7.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X229 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MN1.G xaa6.xf.XA7.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X230 xaa0.xa5.MN0.D xaa0.xa5.MN2.G xaa0.xa5.MP1.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X231 xaa4.xa1.M4.D IBPSR_1U xaa4.xa1.M3.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X232 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R59 xaa4.xa2.M0.G m3_22692_53956# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X233 xaa4.xa1.M8.D xaa1.xa3.D xaa4.xa4.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X234 xaa6.xe.XA6.MN0.G xaa6.xe.XA5.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R60 AVSS m3_37748_88924# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X235 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MN1.G xaa6.xd.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R61 m3_4628_70524# xaa1.xa3.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X236 xaa6.xf.XA7.MN0.D xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X237 xaa5.xa3.xb1_0.G xaa5.xa3.xb2_0.G xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X238 AVDD PWRUP_1V8 xaa6.xe.XA7.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X239 xaa6.xd.XA3.MP0.D xaa6.xd.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X240 xaa3.xa1c.MN0.D xaa3.xa1b.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X241 xaa5.xb2_0.MN0.D xaa5.xb1.MN1.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R62 m3_4628_91644# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X242 a_n508_74698# xbb0.xa1.XA1.N AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X243 xaa6.xe.XA5.MN0.G xaa6.xe.XA7.MN1.G xaa6.xe.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X244 xaa6.xd.XA6.MP0.D xaa6.xd.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X245 xaa5.xa3.xb2_0.G xaa5.xb2_4.MN0.D xaa4.xa2.M0.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X246 xaa5.xa3.xb1_0.D xaa5.xa3.xb1_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X247 xaa3.xa6.MN0.D xaa3.xa1c.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X248 xaa0.xa5.MN2.G xaa6.xc.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X249 AVSS xaa1.xa4.M0.G xaa1.xa4.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X250 xaa6.xc.XA6.MN0.G xaa6.xc.XA5.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R63 AVSS m3_37748_75484# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X251 xaa1.xa2.M1.D IBPSR_1U xaa1.xa2.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X252 xbb1.xa3.M4.D IBPSR_1U xbb1.xa3.M3.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X253 xaa6.xc.XA7.MN1.G PWRUP_1V8 xaa6.xc.XA1.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X254 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X255 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X256 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X257 xaa1.xa1.M8.D xaa1.xa1.M8.D xaa1.xb1.M0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X258 xaa3.xa7.MN0.D xaa3.xa6.MN0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X259 xaa6.xc.XA5.MN0.G xaa6.xc.XA7.MP1.G xaa6.xc.XA4.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R64 m3_4628_83004# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X260 xaa1.xa2.M3.D IBPSR_1U xaa1.xa2.M2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R65 AVSS m3_37748_70684# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X261 xaa1.xa1.M1.D IBPSR_1U xaa1.xa1.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R66 xaa4.xa2.M0.G m3_22692_58180# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X262 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X263 xaa6.xd.XA7.MP1.G xaa6.xd.XA7.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X264 xaa4.xa1.M8.D xaa4.xa2.M0.G xaa4.xa2.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R67 m3_4628_86844# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X265 xaa6.xf.XA6.MN0.G xaa6.xf.XA5.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R68 li_4836_56708# xaa3.xa1c.MN0.D sky130_fd_pr__res_generic_l1 w=0.44 l=0.36
X266 AVDD PWRUP_1V8 xaa6.xf.XA7.MN1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X267 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X268 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
X269 a_1220_70022# a_788_72222# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X270 xaa3.xa9.MN0.D xaa1.xa4.M0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X271 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X272 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MP1.G xaa6.xd.XA6.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X273 xaa6.xg.XA7.MN2.D PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X274 xaa5.xa3.xb1_0.G xaa5.xa3.xb2_0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X275 xaa0.xa6.MN0.D xaa0.xa3.MN1.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X276 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X277 xaa6.xf.XA5.MN0.G xaa6.xf.XA7.MN1.G xaa6.xf.XA4.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X278 xaa6.xe.XA1.MN0.D xaa6.xe.XA1.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X279 xaa6.xd.XA3.MN0.D xaa6.xd.XA7.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X280 xaa6.xg.XA5.MN0.G xaa6.xg.XA3.MN1.G xaa6.xg.XA3.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X281 xaa4.xa4.M0.D xaa1.xa3.D xaa4.xa1.M8.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.616 ps=3.3 w=1.08 l=0.18
X282 a_1220_74698# a_1652_76898# AVSS sky130_fd_pr__res_high_po w=0.72 l=8.8
X283 xaa5.xb2_0.MN0.D xaa5.xb1.MN1.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X284 xaa0.xa2a.MN0.D xaa0.xa2a.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X285 AVDD PWRUP_1V8 xaa6.xc.XA7.MN0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X286 xaa4.xa1.M1.D IBPSR_1U xaa4.xa1.M0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X287 xaa6.xc.XA5.MN0.G xaa6.xc.XA7.MP1.G xaa6.xc.XA3.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X288 xaa5.xa3.xb2_0.D xaa5.xa3.xb1_0.D xaa5.xa3.xc2a.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X289 xaa6.xd.XA6.MN0.D xaa6.xd.XA6.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R69 xaa4.xa2.M0.G m3_22692_55012# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
X290 xaa5.xa3.xb2_0.G xaa5.xb2_4.MN0.D AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X291 xaa1.xa3.D xaa0.xa2a.MN0.D xaa1.xb2.M7.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X292 xaa6.xg.XA7.MP1.G xaa6.xg.XA3.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X293 xaa4.xa2.M0.G xaa4.xa4.M0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
R70 AVSS m3_37748_91804# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X294 xaa6.xg.XA4.MN0.D xaa6.xg.XA4.MN0.G AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R71 m3_4628_78204# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X295 xaa0.xa1.MN0.G xaa0.xa1.MN2.S AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R72 AVSS m3_37748_83164# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X296 xaa6.xc.XA4.MP0.D xaa6.xc.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X297 xaa1.xa1.M6.D IBPSR_1U xaa1.xa1.M5.D AVSS sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X298 xaa5.xa4.MN0.D xaa5.xa3.xb1_0.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X299 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MN1.G xaa6.xg.XA6.MP0.D AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X300 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MN1.G xaa6.xe.XA7.MN0.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X301 xaa1.xa3.D PWRUP_1V8 AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X302 xaa6.xg.XA3.MP0.D xaa6.xg.XA7.MN1.D AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X303 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X304 xaa0.xa6.MN0.D xaa0.xa3.MN1.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X305 xaa1.xa3.D xaa0.xa6.MN0.D xaa1.xa2.M8.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X306 xaa6.xg.XA6.MP0.D xaa6.xg.XA6.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X307 xaa6.xe.XA7.MN0.D xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN2.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
X308 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.616 ps=3.3 w=1.08 l=0.18
X309 xaa0.xa2a.MN0.D xaa0.xa2a.MN0.G AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
R73 m3_4628_73404# xaa1.xa4.M0.D sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
X310 xaa1.xa1.M8.D IBPSR_1U xaa1.xa1.M7.D AVSS sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
C0 AVDD xaa6.xe.XA7.MN1.D 1.86f
C1 CK PWRUP_1V8 0.31f
C2 AVDD a_28612_54510# 0.363f
C3 xaa6.xc.XA7.MN1.G xaa6.xd.XA7.MN1.G 0.31f
C4 xaa6.xg.XA3.MN1.G a_37324_53806# 0.107f
C5 AVDD xaa5.xb1.MN1.D 0.636f
C6 AVDD a_27244_55566# 0.383f
C7 xaa4.xa4.M0.D xaa4.xa2.M0.D 1.3f
C8 AVDD a_28612_56622# 0.365f
C9 AVDD xaa6.xd.XA1.MN0.G 1.64f
C10 AVDD a_27244_54510# 0.363f
C11 xaa6.xc.XA7.MP1.G xaa6.xc.XA7.MN0.D 0.117f
C12 xaa6.xg.XA3.MN1.G a_36172_53806# 0.113f
C13 xaa5.xa3.xb2_0.G a_29764_63566# 0.134f
C14 AVDD PWRUP_1V8 15.3f
C15 AVDD a_27244_56622# 0.365f
C16 AVDD xaa6.xd.XA7.MN1.D 1.86f
C17 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MN0.D 0.336f
C18 xaa4.xa2.M0.G xaa5.xb2_4.MN0.D 0.173f
C19 AVDD xaa6.xg.XA5.MN0.G 0.879f
C20 AVDD a_28612_53102# 0.488f
C21 xaa4.xa4.M0.D a_11784_61708# 0.128f
C22 xaa5.xa3.xb1_0.D a_27244_62158# 0.14f
C23 AVDD xaa6.xc.XA1.MN0.G 3.51f
C24 AVDD xaa6.xg.XA3.MP0.D 0.133f
C25 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MP1.G 0.314f
C26 xaa6.xc.XA7.MN1.G xaa6.xc.XA7.MP1.G 0.537f
C27 AVDD xaa1.xa1.M8.D 2.27f
C28 AVDD xaa6.xg.XA5.MN0.D 0.216f
C29 xaa1.xa4.M0.D m3_37748_87964# 0.111f
C30 AVDD xaa4.xa2.M0.D 5.68f
C31 AVDD a_27244_53102# 0.486f
C32 xaa4.xa2.M0.G m3_13116_55188# 0.106f
C33 AVDD xaa6.xc.XA7.MN1.D 1.86f
C34 xaa6.xg.XA7.MN1.D xaa6.xg.XA7.MN1.G 0.311f
C35 AVDD a_640_61510# 0.333f
C36 AVDD xaa6.xf.XA5.MN0.G 0.88f
C37 a_1652_76898# xaa1.xa4.M0.D 0.163f
C38 AVDD a_37324_56974# 0.405f
C39 xaa0.xa2a.MN0.D xaa0.xa2a.MN0.G 0.14f
C40 IBPSR_1U xaa0.xa2a.MN0.D 0.58f
C41 AVDD xaa0.xa5.MN2.G 4.18f
C42 AVDD xaa6.xg.XA3.MN1.G 1.14f
C43 xaa6.xf.XA1.MN0.G xaa6.xg.XA7.MN1.G 0.128f
C44 AVDD xaa6.xe.XA5.MN0.G 0.88f
C45 AVDD a_37324_58030# 0.344f
C46 xaa6.xc.XA6.MN0.G xaa6.xc.XA5.MN0.G 0.27f
C47 AVDD a_11784_61708# 0.517f
C48 AVDD xaa6.xd.XA5.MN0.G 0.88f
C49 AVDD xaa6.xf.XA3.MP0.D 0.133f
C50 xaa6.xf.XA1.MN0.G xaa6.xf.XA7.MN1.G 0.224f
C51 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MN0.D 0.336f
C52 xaa6.xf.XA6.MN0.G a_33652_55918# 0.111f
C53 xaa1.xa4.M0.D m3_37748_88924# 0.111f
C54 AVDD a_33652_56974# 0.405f
C55 AVDD a_11784_53260# 0.519f
C56 xaa4.xa2.M0.G m3_13116_56244# 0.106f
C57 xaa5.xa3.xb2_0.D xaa5.xa3.xc2a.D 0.123f
C58 AVDD xaa6.xe.XA3.MP0.D 0.133f
C59 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN0.D 0.129f
C60 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MN1.G 0.467f
C61 xaa4.xa2.M0.G xaa5.xa3.xb2_0.G 0.416f
C62 xaa1.xa4.M0.G xaa0.xa6.MN0.D 0.25f
C63 AVDD a_28612_61806# 0.352f
C64 AVDD a_5844_55150# 0.443f
C65 PWRUP_1V8 xaa6.xg.XA7.MP1.G 0.124f
C66 AVDD a_32284_56974# 0.405f
C67 xaa4.xa2.M0.D a_11784_53788# 0.111f
C68 AVDD a_33652_58030# 0.338f
C69 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN1.G 0.201f
C70 xaa6.xf.XA7.MN1.D xaa6.xf.XA7.MP1.G 0.313f
C71 xaa6.xe.XA6.MN0.G a_32284_55918# 0.113f
C72 xaa5.xa3.xb1_0.G xaa5.xa3.xb2_0.G 1.05f
C73 AVDD a_27244_61806# 0.364f
C74 PWRUP_1V8 xaa6.xg.XA7.MN1.G 0.275f
C75 xaa6.xg.XA7.MP1.G xaa6.xg.XA5.MN0.G 0.397f
C76 xbb0.xa1.XA1.N a_n76_72222# 0.113f
C77 AVDD a_32284_58030# 0.343f
C78 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MP1.G 0.216f
C79 xaa1.xa4.M0.D m3_37748_72604# 0.111f
C80 xaa5.xa3.xb1_0.G a_29764_63918# 0.133f
C81 AVDD a_5844_55502# 0.485f
C82 AVDD a_37324_53454# 0.369f
C83 xaa0.xa6.MN0.D xaa0.xa2a.MN0.D 3.25f
C84 AVDD xaa6.xd.XA3.MP0.D 0.133f
C85 AVDD xaa5.xb2_0.MN0.D 0.55f
C86 PWRUP_1V8 xaa6.xf.XA7.MN1.G 0.667f
C87 xaa1.xa4.M0.D m3_37748_89884# 0.111f
C88 AVDD a_28612_56974# 0.405f
C89 xaa1.xa1.M8.D a_640_60278# 0.182f
C90 xaa4.xa2.M0.G m3_13116_57300# 0.106f
C91 xaa5.xa3.xb1_0.G a_26092_61102# 0.173f
C92 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MN0.D 0.336f
C93 AVDD xaa6.xc.XA3.MP0.D 0.133f
C94 xaa6.xg.XA7.MP1.G xaa6.xg.XA3.MN1.G 0.352f
C95 xaa5.xa3.xb1_0.G xaa4.xa2.M0.G 0.414f
C96 AVDD xaa5.xa3.xc2a.D 0.159f
C97 PWRUP_1V8 xaa6.xf.XA7.MP1.G 0.124f
C98 AVDD xaa6.xc.XA5.MN0.G 0.88f
C99 xaa3.xa6.MN0.D xaa3.xa1c.MN0.D 0.187f
C100 a_788_76898# a_1652_76898# 0.107f
C101 AVDD a_27244_56974# 0.405f
C102 xaa4.xa4.M0.D a_11784_58012# 0.128f
C103 AVDD a_28612_58030# 0.338f
C104 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN0.D 0.12f
C105 xaa6.xe.XA1.MN0.G xaa6.xe.XA7.MN1.G 0.412f
C106 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MP1.G 0.313f
C107 xaa6.xg.XA7.MN1.G xaa6.xg.XA3.MN1.G 0.129f
C108 xaa6.xd.XA6.MN0.G a_28612_55918# 0.111f
C109 AVDD a_37324_55918# 0.386f
C110 xaa4.xa4.M0.D a_11784_58540# 0.128f
C111 AVDD a_33652_53454# 0.368f
C112 xaa5.xb2_2.MN0.D xaa5.xb2_1.MN0.D 0.197f
C113 AVDD a_27244_58030# 0.343f
C114 IBPSR_1U PWRUP_1V8 2.41f
C115 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MP1.G 0.21f
C116 xaa6.xe.XA7.MN1.D xaa6.xe.XA7.MN1.G 0.467f
C117 xaa1.xa4.M0.D m3_37748_73564# 0.111f
C118 xaa5.xb1.MN1.G xaa4.xa2.M0.G 0.132f
C119 PWRUP_1V8 xaa6.xe.XA7.MP1.G 0.124f
C120 xaa3.xa6.MN0.D a_4692_58142# 0.117f
C121 AVDD a_11784_56956# 0.517f
C122 xaa4.xa4.M0.D a_11784_59068# 0.128f
C123 AVDD a_32284_53454# 0.367f
C124 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN1.G 0.195f
C125 AVDD a_37324_54862# 0.382f
C126 xaa6.xc.XA6.MN0.G a_27244_55918# 0.113f
C127 xaa5.xb1.MN1.G xaa5.xa3.xb1_0.G 0.194f
C128 AVDD a_28612_62158# 0.352f
C129 PWRUP_1V8 xaa6.xe.XA7.MN1.G 0.658f
C130 xaa3.xa1b.MN0.D xaa3.xa1c.MN0.D 0.406f
C131 xaa6.xf.XA7.MP1.G xaa6.xf.XA5.MN0.G 0.397f
C132 xaa1.xa4.M0.D m3_37748_90844# 0.111f
C133 xbb0.xa1.XA1.N xaa1.xa4.M0.D 0.448f
C134 xaa4.xa4.M0.D a_11784_59596# 0.128f
C135 xaa4.xa2.M0.G m3_13116_58356# 0.106f
C136 AVDD a_11784_58012# 0.517f
C137 PWRUP_1V8 xaa0.xa1.MN0.G 0.238f
C138 AVDD a_27244_62158# 0.384f
C139 AVDD a_33652_55918# 0.385f
C140 a_n940_74698# xaa1.xa4.M0.D 0.187f
C141 AVDD xaa6.xg.XA7.MN0.G 0.479f
C142 xaa0.xa3.MN1.G xaa0.xa5.MN2.D 0.152f
C143 AVDD a_11784_58540# 0.517f
C144 xaa5.xa3.xb2_0.D xaa5.xa3.xb1_0.D 0.607f
C145 xaa4.xa4.M0.D a_11784_62236# 0.128f
C146 xaa6.xd.XA1.MN0.G xaa6.xd.XA7.MN1.G 0.224f
C147 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MN0.D 0.336f
C148 AVDD a_32284_55918# 0.385f
C149 PWRUP_1V8 xaa6.xd.XA7.MN1.G 0.667f
C150 AVDD xaa1.xa4.M0.D 0.873f
C151 AVDD a_28612_53454# 0.368f
C152 xaa0.xa3.MN1.G xaa0.xa5.MN0.D 0.446f
C153 AVDD a_11784_59068# 0.517f
C154 IBPSR_1U a_n908_61510# 0.156f
C155 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN0.D 0.129f
C156 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MN1.G 0.467f
C157 AVDD a_33652_54862# 0.383f
C158 xaa1.xa4.M0.D m3_37748_74524# 0.111f
C159 xaa3.xa1b.MN0.D xaa3.xa6.MN0.D 0.137f
C160 PWRUP_1V8 xaa6.xd.XA7.MP1.G 0.124f
C161 xaa6.xe.XA7.MP1.G xaa6.xe.XA5.MN0.G 0.397f
C162 AVDD a_27244_53454# 0.367f
C163 xaa6.xg.XA5.MN0.G xaa6.xg.XA4.MN0.D 0.126f
C164 AVDD a_11784_59596# 0.517f
C165 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN1.G 0.201f
C166 xaa6.xd.XA7.MN1.D xaa6.xd.XA7.MP1.G 0.313f
C167 xaa6.xg.XA7.MN1.D a_36172_57678# 0.132f
C168 AVDD a_32284_54862# 0.383f
C169 AVDD xaa5.xb2_1.MN0.D 0.543f
C170 xaa1.xa4.M0.D m3_37748_91804# 0.111f
C171 xaa4.xa2.M0.G m3_13116_59412# 0.106f
C172 xaa0.xa6.MN0.D PWRUP_1V8 0.181f
C173 AVDD a_5844_57790# 0.364f
C174 xaa5.xb2_2.MN0.D a_29764_62510# 0.126f
C175 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MP1.G 0.216f
C176 AVDD a_11784_62236# 0.517f
C177 PWRUP_1V8 xaa6.xc.XA7.MP1.G 0.124f
C178 AVDD a_28612_55918# 0.385f
C179 a_n76_76898# a_788_76898# 0.107f
C180 AVDD xaa5.xa3.xb1_0.D 1.88f
C181 PWRUP_1V8 xaa6.xc.XA7.MN1.G 0.671f
C182 AVDD a_27244_55918# 0.385f
C183 AVDD a_244_56270# 0.384f
C184 AVDD xaa3.xa1c.MN0.D 1.12f
C185 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MN0.D 0.336f
C186 AVDD a_28612_54862# 0.383f
C187 xaa6.xf.XA7.MN1.D a_34804_57678# 0.134f
C188 xaa1.xa4.M0.D m3_37748_75484# 0.111f
C189 AVDD xaa5.xa4.MN0.D 0.227f
C190 xaa3.xa7.MN0.D xaa3.xa6.MN0.D 0.128f
C191 xaa6.xf.XA5.MN0.G xaa6.xf.XA4.MN0.D 0.126f
C192 AVDD a_5844_58142# 0.388f
C193 xaa6.xc.XA1.MN0.G xaa6.xc.XA7.MN1.G 0.412f
C194 xaa0.xa5.MN2.G xaa6.xc.XA7.MN0.D 0.12f
C195 AVDD a_27244_54862# 0.383f
C196 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MP1.G 0.313f
C197 xaa1.xa3.D xaa4.xa2.M0.G 0.168f
C198 AVDD a_11784_55900# 0.517f
C199 xaa6.xd.XA7.MP1.G xaa6.xd.XA5.MN0.G 0.397f
C200 xaa1.xa4.M0.D m3_37748_92764# 0.111f
C201 xaa4.xa2.M0.G m3_13116_60468# 0.106f
C202 xaa6.xf.XA7.MN1.G a_33652_53454# 0.101f
C203 xaa4.xa2.M0.G xaa5.xb1.MN1.D 0.226f
C204 xaa0.xa5.MN2.G xaa6.xc.XA7.MP1.G 0.193f
C205 xaa6.xc.XA7.MN1.D xaa6.xc.XA7.MN1.G 0.467f
C206 AVDD xaa6.xg.XA6.MN0.G 0.478f
C207 AVDD xaa0.xa5.MN0.D 0.697f
C208 AVDD xaa3.xa6.MN0.D 0.724f
C209 AVDD a_11784_54844# 0.517f
C210 AVDD xaa6.xf.XA6.MN0.G 1.7f
C211 xaa3.xa7.MN0.D xaa3.xa1b.MN0.D 0.123f
C212 xaa5.xb1.MN1.D xaa5.xb1.MN0.D 0.106f
C213 AVDD a_244_56622# 0.388f
C214 AVDD a_5844_58494# 0.388f
C215 AVDD xaa6.xg.XA4.MN0.G 0.485f
C216 xaa1.xa4.M0.D m3_37748_76444# 0.111f
C217 AVDD a_28612_62510# 0.352f
C218 AVDD xaa6.xe.XA6.MN0.G 1.7f
C219 xaa6.xe.XA5.MN0.G xaa6.xe.XA4.MN0.D 0.126f
C220 xaa5.xb1.MN1.G xaa5.xb1.MN1.D 0.209f
C221 xaa6.xe.XA7.MN1.D a_31132_57678# 0.132f
C222 AVDD a_27244_62510# 0.388f
C223 AVDD xaa6.xd.XA6.MN0.G 1.7f
C224 xaa4.xa2.M0.G xaa4.xa2.M0.D 0.544f
C225 xbb0.xa1.XA1.N a_n76_76898# 0.119f
C226 AVDD xaa0.xa3.MN1.G 1.25f
C227 xaa4.xa2.M0.G m3_13116_61524# 0.106f
C228 AVDD xaa3.xa1b.MN0.D 1.37f
C229 AVDD a_37324_55214# 0.364f
C230 AVDD xaa6.xc.XA6.MN0.G 1.7f
C231 xbb0.xa1.XA1.N a_n508_74698# 0.207f
C232 AVDD a_244_56974# 0.349f
C233 xaa6.xe.XA7.MN1.G a_32284_53454# 0.101f
C234 xaa6.xd.XA5.MN0.G xaa6.xd.XA4.MN0.D 0.126f
C235 AVDD a_5844_58846# 0.364f
C236 xaa6.xf.XA1.MN0.G xaa6.xg.XA7.MN1.D 0.147f
C237 AVDD xaa5.xb2_2.MN0.D 0.543f
C238 AVDD a_37324_56270# 0.362f
C239 PWRUP_1V8 xaa0.xa2a.MN0.D 0.579f
C240 AVDD a_37324_53806# 0.405f
C241 xaa6.xd.XA7.MN1.D a_29764_57678# 0.134f
C242 xaa1.xa4.M0.D m3_37748_77404# 0.111f
C243 xaa4.xa2.M0.D a_11784_55372# 0.138f
C244 AVDD xaa5.xa3.xb2_0.D 1.82f
C245 AVDD a_37324_57326# 0.364f
C246 xaa4.xa2.M0.D a_11784_54316# 0.112f
C247 AVDD xaa3.xa8.MP0.D 0.191f
C248 xaa5.xa3.xb2_0.G a_26092_61806# 0.175f
C249 AVDD a_33652_55214# 0.364f
C250 xaa4.xa2.M0.D xaa4.xa1.M8.D 0.21f
C251 AVDD xaa4.xa4.M0.D 8.82f
C252 xaa6.xg.XA7.MP1.G xaa6.xg.XA6.MN0.G 0.111f
C253 xaa6.xc.XA7.MP1.G xaa6.xc.XA5.MN0.G 0.397f
C254 a_n940_74698# xbb0.xa1.XA1.N 0.104f
C255 xaa6.xg.XA5.MN0.G a_36172_55566# 0.112f
C256 xaa4.xa2.M0.G m3_13116_62580# 0.106f
C257 xaa6.xf.XA7.MN1.G xaa6.xf.XA1.MN0.D 0.123f
C258 AVDD xaa3.xa7.MN0.D 0.714f
C259 AVDD a_32284_55214# 0.364f
C260 AVDD a_33652_56270# 0.363f
C261 xaa4.xa2.M0.D a_11784_56428# 0.142f
C262 xaa5.xb1.MN1.D a_29764_61454# 0.127f
C263 AVDD a_33652_53806# 0.406f
C264 AVDD a_5844_59198# 0.384f
C265 xaa6.xe.XA1.MN0.G xaa6.xf.XA7.MN1.D 0.274f
C266 xaa6.xg.XA7.MP1.G xaa6.xg.XA4.MN0.G 0.127f
C267 AVDD CK 3.95f
C268 xaa1.xa3.D a_2948_70022# 0.202f
C269 PWRUP_1V8 xaa6.xg.XA7.MN1.D 0.16f
C270 AVDD a_32284_56270# 0.363f
C271 AVDD a_33652_57326# 0.364f
C272 xaa3.xa1b.MN0.D a_4692_55854# 0.124f
C273 AVDD a_32284_53806# 0.406f
C274 xaa6.xd.XA7.MN1.G a_28612_53454# 0.101f
C275 xaa3.xa1c.MN0.D li_6204_57236# 0.118f
C276 xaa1.xa4.M0.D m3_37748_78364# 0.111f
C277 AVDD a_11784_62764# 0.428f
C278 PWRUP_1V8 xaa6.xf.XA1.MN0.G 0.456f
C279 xaa6.xg.XA7.MN1.D xaa6.xg.XA5.MN0.G 0.29f
C280 AVDD a_32284_57326# 0.364f
C281 xaa6.xf.XA5.MN0.G a_34804_55566# 0.113f
C282 AVDD xaa3.xa9.MN0.D 0.176f
C283 xaa4.xa2.M0.G xaa5.xb2_0.MN0.D 0.174f
C284 AVDD a_28612_55214# 0.364f
C285 xaa6.xc.XA7.MN1.D a_26092_57678# 0.132f
C286 PWRUP_1V8 xaa6.xf.XA7.MN1.D 0.161f
C287 xaa6.xf.XA7.MN1.G xaa6.xf.XA6.MN0.G 0.329f
C288 xaa4.xa2.M0.G m3_13116_63636# 0.106f
C289 AVDD a_5844_59550# 0.351f
C290 xaa5.xb2_3.MN0.D xaa5.xb2_2.MN0.D 0.197f
C291 AVDD a_27244_55214# 0.364f
C292 AVDD a_28612_62862# 0.352f
C293 PWRUP_1V8 xaa6.xe.XA1.MN0.G 0.209f
C294 AVDD a_28612_56270# 0.363f
C295 xaa6.xf.XA7.MP1.G xaa6.xf.XA6.MN0.G 0.524f
C296 xaa4.xa4.M0.D a_11784_60124# 0.128f
C297 AVDD a_28612_53806# 0.406f
C298 xaa6.xe.XA7.MN1.G xaa6.xe.XA1.MN0.D 0.123f
C299 xaa6.xd.XA1.MN0.G xaa6.xe.XA7.MN1.D 0.262f
C300 xaa6.xg.XA7.MN1.D xaa6.xg.XA3.MN1.G 0.158f
C301 AVDD a_27244_62862# 0.469f
C302 PWRUP_1V8 xaa6.xe.XA7.MN1.D 0.16f
C303 AVDD a_27244_56270# 0.363f
C304 AVDD a_28612_57326# 0.364f
C305 AVDD a_27244_53806# 0.406f
C306 xaa6.xc.XA5.MN0.G xaa6.xc.XA4.MN0.D 0.126f
C307 AVDD a_640_59750# 0.389f
C308 AVDD CK_REF 0.562f
C309 xaa1.xa4.M0.D m3_37748_79324# 0.111f
C310 PWRUP_1V8 xaa6.xd.XA1.MN0.G 0.537f
C311 xaa6.xf.XA7.MN1.D xaa6.xf.XA5.MN0.G 0.29f
C312 AVDD a_27244_57326# 0.364f
C313 xaa6.xe.XA5.MN0.G a_31132_55566# 0.112f
C314 xaa6.xc.XA7.MN1.G a_27244_53454# 0.101f
C315 AVDD a_244_53806# 0.384f
C316 a_1652_72222# xaa1.xa3.D 0.168f
C317 PWRUP_1V8 xaa6.xd.XA7.MN1.D 0.161f
C318 AVDD a_5844_55854# 0.388f
C319 xaa6.xe.XA7.MP1.G xaa6.xe.XA6.MN0.G 0.524f
C320 xaa0.xa5.MN0.D xaa0.xa1.MN0.G 0.15f
C321 AVDD a_11784_53788# 0.517f
C322 xaa6.xd.XA7.MN1.G xaa6.xd.XA1.MN0.D 0.123f
C323 AVDD a_11784_60124# 0.517f
C324 PWRUP_1V8 xaa6.xc.XA1.MN0.G 0.212f
C325 xaa6.xe.XA7.MN1.G xaa6.xe.XA6.MN0.G 0.329f
C326 IBPSR_1U xaa3.xa1b.MN0.D 0.837f
C327 xaa1.xa1.M8.D PWRUP_1V8 0.25f
C328 AVDD xaa6.xg.XA7.MN0.D 0.485f
C329 xaa6.xd.XA5.MN0.G a_29764_55566# 0.113f
C330 xaa6.xc.XA1.MN0.G xaa6.xd.XA7.MN1.D 0.274f
C331 AVDD xaa5.xb2_3.MN0.D 0.545f
C332 PWRUP_1V8 xaa6.xc.XA7.MN1.D 0.162f
C333 CK xaa6.xg.XA7.MN1.G 0.293f
C334 AVDD a_5844_56206# 0.348f
C335 xaa6.xe.XA7.MN1.D xaa6.xe.XA5.MN0.G 0.29f
C336 AVDD xaa6.xg.XA7.MP1.G 2.06f
C337 xaa4.xa4.M0.D a_11784_60652# 0.128f
C338 xaa6.xf.XA7.MN1.G a_34804_53806# 0.115f
C339 xaa6.xg.XA5.MN0.D xaa6.xg.XA5.MN0.G 0.109f
C340 xaa5.xb2_3.MN0.D a_29764_62862# 0.126f
C341 xaa5.xa3.xb2_0.G xaa5.xa3.xb1_0.D 0.294f
C342 AVDD xaa0.xa1.MN0.D 0.702f
C343 xaa1.xa4.M0.D m3_37748_80284# 0.111f
C344 PWRUP_1V8 xaa0.xa5.MN2.G 5.41f
C345 AVDD m1_37504_55818# 0.427f
C346 xaa6.xf.XA7.MP1.G a_34804_56270# 0.1f
C347 PWRUP_1V8 xaa6.xg.XA3.MN1.G 0.382f
C348 xaa0.xa3.MN1.G xaa0.xa1.MN0.G 0.439f
C349 AVDD xaa6.xg.XA7.MN1.G 1.97f
C350 AVDD a_244_52750# 0.443f
C351 xaa6.xf.XA7.MN1.G a_33652_53806# 0.113f
C352 AVDD a_640_60278# 0.385f
C353 xaa4.xa2.M0.G xaa5.xb2_1.MN0.D 0.174f
C354 AVDD a_244_54158# 0.388f
C355 xaa1.xa4.M0.D xaa1.xa4.M0.G 0.231f
C356 AVDD xaa0.xa1.MN2.S 1.24f
C357 AVDD m1_37504_57930# 0.329f
C358 xaa6.xd.XA7.MN1.G xaa6.xd.XA6.MN0.G 0.329f
C359 AVDD xaa6.xf.XA7.MN0.D 0.486f
C360 AVDD a_28612_63214# 0.352f
C361 AVDD a_244_55214# 0.364f
C362 xaa6.xd.XA7.MN1.D xaa6.xd.XA5.MN0.G 0.29f
C363 xaa6.xd.XA7.MP1.G xaa6.xd.XA6.MN0.G 0.524f
C364 AVDD xaa6.xf.XA7.MN1.G 3.56f
C365 AVDD a_244_53102# 0.485f
C366 xaa6.xc.XA7.MN1.G xaa6.xc.XA1.MN0.D 0.123f
C367 AVDD a_11784_60652# 0.517f
C368 AVDD a_244_54510# 0.388f
C369 xaa0.xa5.MN2.G xaa6.xc.XA7.MN1.D 0.248f
C370 AVDD a_27244_63214# 0.439f
C371 xaa0.xa1.MN0.D CK_REF 0.202f
C372 AVDD xaa6.xf.XA7.MP1.G 2.06f
C373 xaa5.xa3.xb1_0.G xaa5.xa3.xb1_0.D 0.192f
C374 xaa1.xa4.M0.D m3_37748_81244# 0.111f
C375 xaa0.xa6.MN0.D xaa0.xa3.MN1.G 0.142f
C376 AVDD xaa0.xa3.MP0.D 0.191f
C377 AVDD xaa6.xe.XA7.MN0.D 0.485f
C378 AVDD a_244_53454# 0.365f
C379 xaa0.xa1.MN2.S CK_REF 0.104f
C380 AVDD a_28612_60750# 0.336f
C381 AVDD xaa0.xa2a.MN0.G 0.717f
C382 a_788_72222# a_1652_72222# 0.107f
C383 AVDD IBPSR_1U 1.83f
C384 AVDD a_244_55566# 0.383f
C385 xaa6.xc.XA7.MP1.G xaa6.xc.XA6.MN0.G 0.524f
C386 xaa4.xa2.M0.D a_11784_53260# 0.111f
C387 AVDD xaa6.xe.XA7.MP1.G 2.06f
C388 xaa5.xb2_0.MN0.D xaa5.xb1.MN1.D 0.184f
C389 xaa6.xg.XA7.MP1.G xaa6.xg.XA7.MN0.D 0.117f
C390 xaa6.xe.XA7.MN1.G a_32284_53806# 0.115f
C391 AVDD a_27244_60750# 0.367f
C392 AVDD a_244_54862# 0.386f
C393 xaa6.xc.XA7.MN1.G xaa6.xc.XA6.MN0.G 0.329f
C394 AVDD xaa6.xe.XA7.MN1.G 3.52f
C395 AVDD xaa0.xa1.MP1.D 0.191f
C396 xaa6.xe.XA7.MN1.G a_31132_53806# 0.114f
C397 AVDD xaa5.xb2_4.MN0.D 0.541f
C398 AVDD xaa0.xa1.MN0.G 1.23f
C399 xaa6.xg.XA7.MP1.G m1_37504_55818# 0.242f
C400 AVDD xaa6.xd.XA7.MN0.D 0.485f
C401 xaa6.xg.XA7.MN1.G xaa6.xg.XA7.MP1.G 0.141f
C402 xaa6.xc.XA5.MN0.G a_26092_55566# 0.112f
C403 xaa0.xa1.MN2.S xaa0.xa1.MN2.D 0.157f
C404 AVDD xaa6.xg.XA4.MP0.D 0.159f
C405 xaa1.xa4.M0.D m3_37748_82204# 0.111f
C406 AVDD a_244_55918# 0.364f
C407 xaa6.xg.XA7.MP1.G m1_37504_57930# 0.13f
C408 xaa6.xg.XA7.MN1.G m1_37504_55818# 0.153f
C409 AVDD xaa6.xd.XA7.MN1.G 3.56f
C410 AVDD a_37324_54158# 0.386f
C411 xaa1.xa3.D m3_37748_69724# 0.111f
C412 xaa0.xa1.MN2.S xaa0.xa1.MN0.D 0.423f
C413 xaa5.xa3.xb2_0.G xaa5.xa3.xb2_0.D 0.145f
C414 AVDD xaa6.xd.XA7.MP1.G 2.06f
C415 xaa6.xd.XA7.MN1.G a_29764_53806# 0.115f
C416 AVDD xaa6.xg.XA4.MP1.G 0.349f
C417 AVDD a_28612_63566# 0.351f
C418 AVDD xaa0.xa5.MP1.D 0.191f
C419 xaa4.xa4.M0.D a_11784_57484# 0.128f
C420 xaa6.xd.XA7.MP1.G a_29764_56270# 0.1f
C421 xaa6.xc.XA7.MN1.D xaa6.xc.XA5.MN0.G 0.29f
C422 AVDD xaa6.xc.XA7.MN0.D 0.485f
C423 xaa5.xa3.xb2_0.D a_27244_61102# 0.164f
C424 xaa0.xa1.MN0.G CK_REF 0.13f
C425 xaa6.xd.XA7.MN1.G a_28612_53806# 0.113f
C426 AVDD a_640_60806# 0.356f
C427 xaa4.xa2.M0.G xaa5.xb2_2.MN0.D 0.174f
C428 AVDD xaa0.xa6.MN0.D 1.43f
C429 xaa1.xa4.M0.D xaa1.xa3.D 4f
C430 AVDD xaa6.xg.XA6.MP0.D 0.147f
C431 AVDD a_37324_52750# 0.448f
C432 AVDD xaa6.xc.XA7.MP1.G 2.06f
C433 AVDD a_33652_54158# 0.387f
C434 AVDD xaa6.xf.XA4.MP0.D 0.159f
C435 xaa1.xa4.M0.D m3_37748_83164# 0.111f
C436 xaa5.xb2_0.MN0.D a_29764_61806# 0.126f
C437 AVDD xaa6.xc.XA7.MN1.G 3.53f
C438 xaa6.xf.XA7.MP1.G xaa6.xf.XA7.MN0.D 0.117f
C439 AVDD a_32284_54158# 0.387f
C440 xaa1.xa3.D m3_37748_70684# 0.111f
C441 xaa4.xa2.M0.G xaa4.xa4.M0.D 1.94f
C442 AVDD xaa6.xe.XA4.MP0.D 0.159f
C443 AVDD xaa5.xa3.xb2_0.G 0.952f
C444 a_n76_72222# a_788_72222# 0.107f
C445 xaa5.xa3.xb1_0.D a_27244_61454# 0.113f
C446 AVDD a_11784_57484# 0.517f
C447 xaa6.xf.XA7.MP1.G xaa6.xf.XA7.MN1.G 0.537f
C448 xaa0.xa1.MN2.S xaa0.xa2a.MN0.G 0.405f
C449 AVDD a_28612_61102# 0.352f
C450 xaa5.xb2_4.MN0.D xaa5.xb2_3.MN0.D 0.197f
C451 AVDD xaa6.xf.XA6.MP0.D 0.147f
C452 AVDD a_33652_52750# 0.447f
C453 AVDD a_37324_57678# 0.383f
C454 xaa0.xa1.MN0.G xaa0.xa1.MN0.D 0.274f
C455 AVDD a_27244_61102# 0.363f
C456 xaa4.xa2.M0.G CK 0.794f
C457 AVDD a_28612_63918# 0.351f
C458 AVDD xaa6.xe.XA6.MP0.D 0.147f
C459 AVDD a_32284_52750# 0.449f
C460 xaa1.xa4.M0.G xaa3.xa7.MN0.D 0.347f
C461 AVDD a_28612_54158# 0.387f
C462 xaa6.xc.XA7.MN1.G a_27244_53806# 0.115f
C463 xaa5.xa3.xb1_0.G CK 0.129f
C464 xaa5.xb2_4.MN0.D a_29764_63214# 0.126f
C465 AVDD xaa6.xd.XA4.MP0.D 0.159f
C466 xaa1.xa4.M0.D m3_37748_84124# 0.111f
C467 AVDD xaa4.xa2.M0.G 11f
C468 xaa0.xa2a.MN0.G a_n908_54510# 0.112f
C469 xaa4.xa4.M0.D a_11784_61180# 0.128f
C470 xaa6.xe.XA7.MN1.G xaa6.xf.XA7.MN1.G 0.31f
C471 xaa4.xa4.M0.D xaa4.xa1.M8.D 0.217f
C472 AVDD a_27244_54158# 0.387f
C473 xaa1.xa3.D m3_37748_71644# 0.111f
C474 xaa6.xc.XA7.MN1.G a_26092_53806# 0.114f
C475 AVDD xaa1.xb2.M7.D 0.166f
C476 AVDD xaa6.xc.XA4.MP0.D 0.159f
C477 AVDD xaa5.xa3.xb1_0.G 0.826f
C478 xaa6.xf.XA7.MN1.D xaa6.xf.XA6.MN0.G 0.224f
C479 AVDD a_33652_57678# 0.384f
C480 xaa6.xe.XA7.MP1.G xaa6.xe.XA7.MN0.D 0.117f
C481 AVDD xaa1.xa4.M0.G 2.39f
C482 AVDD xaa6.xd.XA6.MP0.D 0.147f
C483 AVDD a_28612_52750# 0.447f
C484 AVDD a_32284_57678# 0.384f
C485 xaa1.xa4.M0.G xaa3.xa9.MN0.D 0.169f
C486 AVDD xaa5.xa3.xc1a.D 0.153f
C487 AVDD a_11784_55372# 0.517f
C488 AVDD xaa5.xb1.MN1.G 0.635f
C489 AVDD xaa6.xc.XA6.MP0.D 0.147f
C490 AVDD a_27244_52750# 0.449f
C491 AVDD a_11784_54316# 0.517f
C492 xaa6.xe.XA7.MN1.G xaa6.xe.XA7.MP1.G 0.537f
C493 xaa6.xg.XA3.MN1.G xaa6.xg.XA1.MN0.D 0.122f
C494 AVDD a_11784_61180# 0.517f
C495 xaa1.xa4.M0.D m3_37748_85084# 0.111f
C496 IBPSR_1U a_4308_51918# 0.136f
C497 xaa6.xe.XA7.MN1.D xaa6.xe.XA6.MN0.G 0.224f
C498 AVDD xaa0.xa2a.MN0.D 1.72f
C499 AVDD a_37324_55566# 0.383f
C500 xaa4.xa2.M0.D a_11784_55900# 0.142f
C501 AVDD a_11784_56428# 0.517f
C502 AVDD a_11784_52732# 0.497f
C503 AVDD a_28612_57678# 0.384f
C504 AVDD a_37324_54510# 0.362f
C505 AVDD a_28612_64270# 0.351f
C506 AVDD a_37324_56622# 0.364f
C507 AVDD a_27244_57678# 0.384f
C508 xaa4.xa2.M0.D a_11784_54844# 0.12f
C509 xaa4.xa2.M0.G xaa5.xb2_3.MN0.D 0.174f
C510 AVDD a_640_61158# 0.376f
C511 AVDD xaa5.xb3.MP1.D 0.476f
C512 PWRUP_1V8 xaa3.xa1b.MN0.D 1.73f
C513 xaa6.xd.XA7.MN1.D xaa6.xd.XA6.MN0.G 0.224f
C514 xaa0.xa5.MN2.G xaa0.xa5.MN0.D 0.22f
C515 xaa6.xf.XA6.MN0.G xaa6.xf.XA5.MN0.G 0.27f
C516 xaa0.xa6.MN0.D IBPSR_1U 0.226f
C517 AVDD a_33652_55566# 0.383f
C518 xaa1.xa4.M0.D m3_37748_86044# 0.111f
C519 AVDD a_37324_53102# 0.485f
C520 xaa4.xa2.M0.G m3_13116_53076# 0.106f
C521 xaa5.xb2_1.MN0.D xaa5.xb2_0.MN0.D 0.197f
C522 AVDD xaa6.xg.XA7.MN1.D 1.86f
C523 xaa5.xa3.xb1_0.D a_27244_61806# 0.154f
C524 AVDD a_33652_54510# 0.363f
C525 xaa6.xd.XA7.MP1.G xaa6.xd.XA7.MN0.D 0.117f
C526 AVDD a_32284_55566# 0.383f
C527 AVDD a_28612_64622# 0.335f
C528 AVDD a_33652_56622# 0.365f
C529 AVDD xaa6.xf.XA1.MN0.G 0.757f
C530 AVDD a_32284_54510# 0.363f
C531 xaa6.xd.XA7.MP1.G xaa6.xd.XA7.MN1.G 0.537f
C532 xaa6.xe.XA6.MN0.G xaa6.xe.XA5.MN0.G 0.27f
C533 AVDD a_28612_61454# 0.352f
C534 xaa1.xa4.M0.D a_n940_70022# 0.181f
C535 AVDD a_32284_56622# 0.365f
C536 xaa6.xc.XA7.MN1.D xaa6.xc.XA6.MN0.G 0.224f
C537 AVDD xaa6.xf.XA7.MN1.D 1.86f
C538 xaa0.xa5.MN2.G xaa0.xa3.MN1.G 0.116f
C539 AVDD a_27244_61454# 0.382f
C540 xaa1.xa4.M0.D a_2948_74698# 0.383f
C541 AVDD a_33652_53102# 0.488f
C542 AVDD xaa6.xe.XA1.MN0.G 3.52f
C543 xaa5.xb2_1.MN0.D a_29764_62158# 0.126f
C544 xaa6.xd.XA6.MN0.G xaa6.xd.XA5.MN0.G 0.27f
C545 xaa5.xa3.xb2_0.G xaa5.xb2_4.MN0.D 0.228f
C546 AVDD a_28612_55566# 0.383f
C547 xaa1.xa4.M0.D m3_37748_87004# 0.111f
C548 AVDD xaa1.xa3.D 3.13f
C549 AVDD a_32284_53102# 0.486f
C550 xaa4.xa2.M0.G m3_13116_54132# 0.106f
C551 m3_22692_52900# AVSS 0.174f
C552 m3_22692_53956# AVSS 0.174f
C553 m3_22692_55012# AVSS 0.174f
C554 m3_22692_56068# AVSS 0.174f
C555 m3_22692_57124# AVSS 0.174f
C556 m3_22692_58180# AVSS 0.174f
C557 m3_22692_59236# AVSS 0.174f
C558 m3_22692_60292# AVSS 0.174f
C559 m3_22692_61348# AVSS 0.174f
C560 m3_22692_62404# AVSS 0.174f
C561 m3_22692_63460# AVSS 0.174f
C562 m3_4628_69564# AVSS 0.189f
C563 m3_4628_70524# AVSS 0.189f
C564 m3_4628_71484# AVSS 0.189f
C565 m3_4628_72444# AVSS 0.189f
C566 m3_4628_73404# AVSS 0.189f
C567 m3_4628_74364# AVSS 0.189f
C568 m3_4628_75324# AVSS 0.189f
C569 m3_4628_76284# AVSS 0.189f
C570 m3_4628_77244# AVSS 0.189f
C571 m3_4628_78204# AVSS 0.189f
C572 m3_4628_79164# AVSS 0.189f
C573 m3_4628_80124# AVSS 0.189f
C574 m3_4628_81084# AVSS 0.189f
C575 m3_4628_82044# AVSS 0.189f
C576 m3_4628_83004# AVSS 0.189f
C577 m3_4628_83964# AVSS 0.189f
C578 m3_4628_84924# AVSS 0.189f
C579 m3_4628_85884# AVSS 0.189f
C580 m3_4628_86844# AVSS 0.189f
C581 m3_4628_87804# AVSS 0.189f
C582 m3_4628_88764# AVSS 0.189f
C583 m3_4628_89724# AVSS 0.189f
C584 m3_4628_90684# AVSS 0.189f
C585 m3_4628_91644# AVSS 0.189f
C586 m3_4628_92604# AVSS 0.189f
C587 li_4836_56708# AVSS 0.115f
C588 a_4308_51566# AVSS 0.491f $ **FLOATING
C589 a_4308_51918# AVSS 0.389f $ **FLOATING
C590 a_37324_52750# AVSS 0.129f $ **FLOATING
C591 a_36172_52750# AVSS 0.572f $ **FLOATING
C592 a_34804_52750# AVSS 0.573f $ **FLOATING
C593 a_33652_52750# AVSS 0.127f $ **FLOATING
C594 a_32284_52750# AVSS 0.127f $ **FLOATING
C595 a_31132_52750# AVSS 0.572f $ **FLOATING
C596 a_29764_52750# AVSS 0.576f $ **FLOATING
C597 a_28612_52750# AVSS 0.127f $ **FLOATING
C598 a_27244_52750# AVSS 0.127f $ **FLOATING
C599 a_26092_52750# AVSS 0.573f $ **FLOATING
C600 a_11784_52732# AVSS 0.17f $ **FLOATING
C601 a_10092_52750# AVSS 0.514f $ **FLOATING
C602 a_36172_53102# AVSS 0.49f $ **FLOATING
C603 a_34804_53102# AVSS 0.488f $ **FLOATING
C604 a_31132_53102# AVSS 0.49f $ **FLOATING
C605 a_29764_53102# AVSS 0.488f $ **FLOATING
C606 a_26092_53102# AVSS 0.49f $ **FLOATING
C607 a_36172_53454# AVSS 0.365f $ **FLOATING
C608 a_34804_53454# AVSS 0.365f $ **FLOATING
C609 a_31132_53454# AVSS 0.364f $ **FLOATING
C610 a_29764_53454# AVSS 0.365f $ **FLOATING
C611 a_26092_53454# AVSS 0.365f $ **FLOATING
C612 xaa6.xg.XA1.MN0.D AVSS 0.169f
C613 xaa6.xf.XA1.MN0.D AVSS 0.169f
C614 xaa6.xe.XA1.MN0.D AVSS 0.15f
C615 xaa6.xd.XA1.MN0.D AVSS 0.169f
C616 xaa6.xc.XA1.MN0.D AVSS 0.15f
C617 a_36172_53806# AVSS 0.384f $ **FLOATING
C618 a_34804_53806# AVSS 0.384f $ **FLOATING
C619 a_31132_53806# AVSS 0.383f $ **FLOATING
C620 a_29764_53806# AVSS 0.384f $ **FLOATING
C621 a_26092_53806# AVSS 0.383f $ **FLOATING
C622 a_4308_53678# AVSS 0.47f $ **FLOATING
C623 a_244_52750# AVSS 0.13f $ **FLOATING
C624 a_n908_52750# AVSS 0.573f $ **FLOATING
C625 a_n908_53102# AVSS 0.49f $ **FLOATING
C626 a_n908_53454# AVSS 0.363f $ **FLOATING
C627 a_36172_54158# AVSS 0.387f $ **FLOATING
C628 a_34804_54158# AVSS 0.387f $ **FLOATING
C629 a_31132_54158# AVSS 0.387f $ **FLOATING
C630 a_29764_54158# AVSS 0.387f $ **FLOATING
C631 a_26092_54158# AVSS 0.388f $ **FLOATING
C632 a_36172_54510# AVSS 0.364f $ **FLOATING
C633 a_34804_54510# AVSS 0.364f $ **FLOATING
C634 a_31132_54510# AVSS 0.364f $ **FLOATING
C635 a_29764_54510# AVSS 0.364f $ **FLOATING
C636 a_26092_54510# AVSS 0.365f $ **FLOATING
C637 xaa6.xg.XA3.MN0.D AVSS 0.162f
C638 xaa6.xg.XA3.MN1.G AVSS 1.62f
C639 xaa6.xf.XA3.MN0.D AVSS 0.162f
C640 xaa6.xe.XA3.MN0.D AVSS 0.162f
C641 xaa6.xd.XA3.MN0.D AVSS 0.162f
C642 xaa6.xc.XA3.MN0.D AVSS 0.162f
C643 a_10092_54510# AVSS 0.372f $ **FLOATING
C644 a_36172_54862# AVSS 0.383f $ **FLOATING
C645 a_34804_54862# AVSS 0.383f $ **FLOATING
C646 a_31132_54862# AVSS 0.383f $ **FLOATING
C647 a_29764_54862# AVSS 0.383f $ **FLOATING
C648 a_26092_54862# AVSS 0.384f $ **FLOATING
C649 xaa6.xg.XA4.MN0.G AVSS 0.53f
C650 a_10092_55038# AVSS 0.365f $ **FLOATING
C651 a_36172_55214# AVSS 0.364f $ **FLOATING
C652 a_34804_55214# AVSS 0.364f $ **FLOATING
C653 a_31132_55214# AVSS 0.364f $ **FLOATING
C654 a_29764_55214# AVSS 0.364f $ **FLOATING
C655 a_26092_55214# AVSS 0.364f $ **FLOATING
C656 CK_REF AVSS 0.957f
C657 a_n908_53806# AVSS 0.363f $ **FLOATING
C658 xaa0.xa1.MN2.D AVSS 0.138f
C659 xaa0.xa1.MN0.D AVSS 1.16f
C660 a_n908_54158# AVSS 0.406f $ **FLOATING
C661 a_n908_54510# AVSS 0.386f $ **FLOATING
C662 xaa0.xa2a.MN0.G AVSS 1.03f
C663 a_n908_54862# AVSS 0.384f $ **FLOATING
C664 xaa6.xg.XA4.MN0.D AVSS 0.139f
C665 xaa6.xf.XA4.MN0.D AVSS 0.139f
C666 xaa6.xe.XA4.MN0.D AVSS 0.139f
C667 xaa6.xd.XA4.MN0.D AVSS 0.139f
C668 xaa6.xc.XA4.MN0.D AVSS 0.139f
C669 xaa4.xa1.M8.D AVSS 0.475f
C670 a_36172_55566# AVSS 0.383f $ **FLOATING
C671 a_34804_55566# AVSS 0.383f $ **FLOATING
C672 a_31132_55566# AVSS 0.383f $ **FLOATING
C673 a_29764_55566# AVSS 0.383f $ **FLOATING
C674 a_26092_55566# AVSS 0.383f $ **FLOATING
C675 xaa6.xg.XA5.MN0.G AVSS 1.26f
C676 xaa6.xg.XA5.MN0.D AVSS 0.229f
C677 xaa6.xf.XA5.MN0.G AVSS 1.25f
C678 xaa6.xe.XA5.MN0.G AVSS 1.26f
C679 xaa6.xd.XA5.MN0.G AVSS 1.25f
C680 a_10092_55566# AVSS 0.425f $ **FLOATING
C681 a_5844_55150# AVSS 0.132f $ **FLOATING
C682 a_4692_55150# AVSS 0.57f $ **FLOATING
C683 a_4692_55502# AVSS 0.49f $ **FLOATING
C684 xaa6.xc.XA5.MN0.G AVSS 1.26f
C685 a_36172_55918# AVSS 0.387f $ **FLOATING
C686 a_34804_55918# AVSS 0.387f $ **FLOATING
C687 a_31132_55918# AVSS 0.387f $ **FLOATING
C688 a_29764_55918# AVSS 0.387f $ **FLOATING
C689 a_26092_55918# AVSS 0.388f $ **FLOATING
C690 xaa6.xg.XA6.MN0.G AVSS 0.523f
C691 xaa6.xf.XA6.MN0.G AVSS 1.29f
C692 xaa6.xe.XA6.MN0.G AVSS 1.29f
C693 xaa6.xd.XA6.MN0.G AVSS 1.29f
C694 xaa6.xc.XA6.MN0.G AVSS 1.29f
C695 a_36172_56270# AVSS 0.362f $ **FLOATING
C696 a_34804_56270# AVSS 0.362f $ **FLOATING
C697 a_31132_56270# AVSS 0.362f $ **FLOATING
C698 a_29764_56270# AVSS 0.362f $ **FLOATING
C699 a_26092_56270# AVSS 0.363f $ **FLOATING
C700 a_4692_55854# AVSS 0.386f $ **FLOATING
C701 a_4692_56206# AVSS 0.436f $ **FLOATING
C702 xaa0.xa1.MN2.S AVSS 1.79f
C703 a_n908_55214# AVSS 0.367f $ **FLOATING
C704 a_n908_55566# AVSS 0.407f $ **FLOATING
C705 xaa0.xa1.MN0.G AVSS 2.58f
C706 a_n908_55918# AVSS 0.362f $ **FLOATING
C707 xaa6.xg.XA6.MN0.D AVSS 0.146f
C708 xaa6.xf.XA6.MN0.D AVSS 0.146f
C709 xaa6.xe.XA6.MN0.D AVSS 0.146f
C710 xaa6.xd.XA6.MN0.D AVSS 0.146f
C711 xaa6.xc.XA6.MN0.D AVSS 0.146f
C712 a_36172_56622# AVSS 0.382f $ **FLOATING
C713 a_34804_56622# AVSS 0.382f $ **FLOATING
C714 a_31132_56622# AVSS 0.382f $ **FLOATING
C715 a_29764_56622# AVSS 0.382f $ **FLOATING
C716 a_26092_56622# AVSS 0.382f $ **FLOATING
C717 xaa4.xa2.M0.D AVSS 1.19f
C718 a_36172_56974# AVSS 0.362f $ **FLOATING
C719 a_34804_56974# AVSS 0.362f $ **FLOATING
C720 a_31132_56974# AVSS 0.362f $ **FLOATING
C721 a_29764_56974# AVSS 0.362f $ **FLOATING
C722 a_26092_56974# AVSS 0.363f $ **FLOATING
C723 xaa6.xg.XA7.MN2.D AVSS 0.181f
C724 xaa6.xg.XA7.MN0.G AVSS 0.51f
C725 xaa6.xf.XA7.MN2.D AVSS 0.181f
C726 xaa6.xe.XA7.MN2.D AVSS 0.181f
C727 xaa6.xd.XA7.MN2.D AVSS 0.181f
C728 xaa6.xc.XA7.MN2.D AVSS 0.181f
C729 a_n908_56270# AVSS 0.362f $ **FLOATING
C730 xaa0.xa5.MN2.D AVSS 0.152f
C731 xaa0.xa5.MN0.D AVSS 1.16f
C732 a_n908_56622# AVSS 0.407f $ **FLOATING
C733 xaa0.xa3.MN1.G AVSS 2.02f
C734 a_244_56974# AVSS 0.129f $ **FLOATING
C735 a_n908_56974# AVSS 0.465f $ **FLOATING
C736 a_36172_57326# AVSS 0.359f $ **FLOATING
C737 a_34804_57326# AVSS 0.359f $ **FLOATING
C738 a_31132_57326# AVSS 0.359f $ **FLOATING
C739 a_29764_57326# AVSS 0.359f $ **FLOATING
C740 a_26092_57326# AVSS 0.36f $ **FLOATING
C741 xaa6.xg.XA7.MN0.D AVSS 0.248f
C742 xaa6.xg.XA7.MP1.G AVSS 1.85f
C743 xaa6.xg.XA7.MN1.G AVSS 1.35f
C744 xaa6.xf.XA7.MN0.D AVSS 0.248f
C745 xaa6.xf.XA7.MN1.G AVSS 2.9f
C746 xaa6.xf.XA7.MP1.G AVSS 1.85f
C747 xaa6.xe.XA7.MN0.D AVSS 0.248f
C748 xaa6.xe.XA7.MP1.G AVSS 1.85f
C749 xaa6.xe.XA7.MN1.G AVSS 2.91f
C750 xaa6.xd.XA7.MN0.D AVSS 0.248f
C751 xaa6.xd.XA7.MN1.G AVSS 2.9f
C752 xaa6.xd.XA7.MP1.G AVSS 1.85f
C753 xaa6.xc.XA7.MN0.D AVSS 0.248f
C754 xaa6.xc.XA7.MP1.G AVSS 1.85f
C755 xaa6.xc.XA7.MN1.G AVSS 3.02f
C756 a_36172_57678# AVSS 0.381f $ **FLOATING
C757 a_34804_57678# AVSS 0.381f $ **FLOATING
C758 a_31132_57678# AVSS 0.381f $ **FLOATING
C759 a_29764_57678# AVSS 0.381f $ **FLOATING
C760 a_26092_57678# AVSS 0.382f $ **FLOATING
C761 xaa6.xg.XA7.MN1.D AVSS 2.68f
C762 xaa6.xf.XA1.MN0.G AVSS 2.93f
C763 xaa6.xf.XA7.MN1.D AVSS 2.67f
C764 xaa6.xe.XA1.MN0.G AVSS 2.89f
C765 xaa6.xe.XA7.MN1.D AVSS 2.68f
C766 xaa6.xd.XA1.MN0.G AVSS 3.54f
C767 xaa6.xd.XA7.MN1.D AVSS 2.67f
C768 xaa6.xc.XA1.MN0.G AVSS 3.02f
C769 xaa6.xc.XA7.MN1.D AVSS 2.67f
C770 xaa0.xa5.MN2.G AVSS 15.3f
C771 a_37324_58030# AVSS 0.129f $ **FLOATING
C772 a_36172_58030# AVSS 0.462f $ **FLOATING
C773 a_34804_58030# AVSS 0.463f $ **FLOATING
C774 a_33652_58030# AVSS 0.127f $ **FLOATING
C775 a_32284_58030# AVSS 0.127f $ **FLOATING
C776 a_31132_58030# AVSS 0.462f $ **FLOATING
C777 a_29764_58030# AVSS 0.463f $ **FLOATING
C778 a_28612_58030# AVSS 0.131f $ **FLOATING
C779 a_27244_58030# AVSS 0.127f $ **FLOATING
C780 a_26092_58030# AVSS 0.465f $ **FLOATING
C781 a_5844_57790# AVSS 0.109f $ **FLOATING
C782 a_4692_57790# AVSS 0.472f $ **FLOATING
C783 xaa3.xa1c.MN0.D AVSS 5.24f
C784 a_4692_58142# AVSS 0.385f $ **FLOATING
C785 xaa3.xa6.MN0.D AVSS 1.11f
C786 a_4692_58494# AVSS 0.384f $ **FLOATING
C787 xaa3.xa1b.MN0.D AVSS 5.25f
C788 a_4692_58846# AVSS 0.369f $ **FLOATING
C789 xaa3.xa7.MN0.D AVSS 1.03f
C790 a_4692_59198# AVSS 0.407f $ **FLOATING
C791 xaa3.xa9.MN0.D AVSS 0.29f
C792 a_5844_59550# AVSS 0.129f $ **FLOATING
C793 a_4692_59550# AVSS 0.468f $ **FLOATING
C794 a_640_59750# AVSS 0.13f $ **FLOATING
C795 a_n908_59750# AVSS 0.519f $ **FLOATING
C796 a_29764_60750# AVSS 0.493f $ **FLOATING
C797 a_28612_60750# AVSS 0.136f $ **FLOATING
C798 a_27244_60750# AVSS 0.127f $ **FLOATING
C799 a_26092_60750# AVSS 0.492f $ **FLOATING
C800 a_29764_61102# AVSS 0.366f $ **FLOATING
C801 a_26092_61102# AVSS 0.384f $ **FLOATING
C802 xaa5.xb1.MN0.D AVSS 0.175f
C803 xaa0.xa2a.MN0.D AVSS 3.65f
C804 a_29764_61454# AVSS 0.38f $ **FLOATING
C805 a_26092_61454# AVSS 0.389f $ **FLOATING
C806 xaa5.xb1.MN1.D AVSS 0.983f
C807 PWRUP_1V8 AVSS 37f
C808 xaa1.xa1.M8.D AVSS 0.735f
C809 a_n908_61510# AVSS 0.398f $ **FLOATING
C810 a_29764_61806# AVSS 0.384f $ **FLOATING
C811 a_26092_61806# AVSS 0.388f $ **FLOATING
C812 xaa5.xb2_0.MN0.D AVSS 0.897f
C813 a_29764_62158# AVSS 0.384f $ **FLOATING
C814 a_26092_62158# AVSS 0.384f $ **FLOATING
C815 xaa5.xb2_1.MN0.D AVSS 0.893f
C816 xaa5.xa3.xb1_0.D AVSS 1.91f
C817 xaa5.xa4.MN0.D AVSS 0.216f
C818 a_29764_62510# AVSS 0.384f $ **FLOATING
C819 a_26092_62510# AVSS 0.388f $ **FLOATING
C820 xaa5.xb2_2.MN0.D AVSS 0.893f
C821 xaa5.xa3.xb2_0.D AVSS 1.43f
C822 xaa4.xa4.M0.D AVSS 1.74f
C823 CK AVSS 13.3f
C824 a_11784_62764# AVSS 0.106f $ **FLOATING
C825 a_29764_62862# AVSS 0.384f $ **FLOATING
C826 a_26092_62862# AVSS 0.467f $ **FLOATING
C827 xaa5.xb2_3.MN0.D AVSS 0.893f
C828 a_29764_63214# AVSS 0.384f $ **FLOATING
C829 a_26092_63214# AVSS 0.531f $ **FLOATING
C830 IBPSR_1U AVSS 23.7f
C831 a_n908_63270# AVSS 0.367f $ **FLOATING
C832 xaa5.xb2_4.MN0.D AVSS 0.893f
C833 xaa1.xa2.M8.D AVSS 0.166f
C834 a_29764_63566# AVSS 0.381f $ **FLOATING
C835 xaa0.xa6.MN0.D AVSS 3.79f
C836 a_n908_63622# AVSS 0.384f $ **FLOATING
C837 xaa5.xa3.xb2_0.G AVSS 3.22f
C838 a_29764_63918# AVSS 0.381f $ **FLOATING
C839 xaa4.xa2.M0.G AVSS 0.958p
C840 xaa5.xa3.xb1_0.G AVSS 3.71f
C841 xaa1.xa4.M0.G AVSS 7.93f
C842 xaa5.xb1.MN1.G AVSS 2.59f
C843 a_n908_64150# AVSS 0.487f $ **FLOATING
C844 a_29764_64270# AVSS 0.469f $ **FLOATING
C845 xaa5.xb3.MP1.D AVSS 0.119f
C846 a_29764_64622# AVSS 0.568f $ **FLOATING
C847 a_28612_64622# AVSS 0.128f $ **FLOATING
C848 a_2948_70022# AVSS 2.6f $ **FLOATING
C849 xaa1.xa3.D AVSS 0.931p
C850 a_2084_70022# AVSS 0.843f
C851 a_1652_72222# AVSS 1.08f
C852 a_1220_70022# AVSS 0.778f
C853 a_788_72222# AVSS 1.08f
C854 a_356_70022# AVSS 0.778f
C855 a_n76_72222# AVSS 1.08f
C856 a_n508_70022# AVSS 0.843f
C857 a_n940_70022# AVSS 2.59f $ **FLOATING
C858 a_2948_74698# AVSS 2.6f $ **FLOATING
C859 xaa1.xa4.M0.D AVSS 6.7p
C860 a_2084_74698# AVSS 0.843f
C861 a_1652_76898# AVSS 1.08f
C862 a_1220_74698# AVSS 0.778f
C863 a_788_76898# AVSS 1.08f
C864 a_356_74698# AVSS 0.778f
C865 a_n76_76898# AVSS 1.08f
C866 a_n508_74698# AVSS 0.843f
C867 xbb0.xa1.XA1.N AVSS 3.4f
C868 a_n940_74698# AVSS 2.59f $ **FLOATING
C869 AVDD AVSS 0.413p
.ends

