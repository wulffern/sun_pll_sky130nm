magic
tech sky130B
magscale 1 1
timestamp 1720908000
<< checkpaint >>
rect 0 0 20276 12444
<< locali >>
rect 20126 0 20276 12444
rect 0 0 20276 150
rect 0 12294 20276 12444
rect 0 0 150 12444
rect 20126 0 20276 12444
rect 150 230 230 286
rect 150 2568 230 2624
rect 2258 4279 2546 4389
rect 2258 1941 2546 2051
<< m3 >>
rect 11560 0 11668 242
rect 19994 202 20164 240
rect 19994 682 20164 720
rect 19994 1162 20164 1200
rect 19994 1642 20164 1680
rect 19994 2122 20164 2160
rect 19994 2602 20164 2640
rect 19994 3082 20164 3120
rect 19994 3562 20164 3600
rect 19994 4042 20164 4080
rect 19994 4522 20164 4560
rect 19994 5002 20164 5040
rect 19994 5482 20164 5520
rect 19994 5962 20164 6000
rect 19994 6442 20164 6480
rect 19994 6922 20164 6960
rect 19994 7402 20164 7440
rect 19994 7882 20164 7920
rect 19994 8362 20164 8400
rect 19994 8842 20164 8880
rect 19994 9322 20164 9360
rect 19994 9802 20164 9840
rect 19994 10282 20164 10320
rect 19994 10762 20164 10800
rect 19994 11242 20164 11280
rect 19994 11722 20164 11760
<< m1 >>
rect 576 1941 754 1971
rect 576 4279 754 4309
rect 754 1941 784 4309
rect 2304 4279 2380 4309
rect 2380 2042 3284 2072
rect 2380 2522 3284 2552
rect 2380 3002 3284 3032
rect 2380 3482 3284 3512
rect 2380 3962 3284 3992
rect 2380 4442 3284 4472
rect 2380 4922 3284 4952
rect 2380 5402 3284 5432
rect 2380 5882 3284 5912
rect 2380 6362 3284 6392
rect 2380 6842 3284 6872
rect 2380 7322 3284 7352
rect 2380 7802 3284 7832
rect 2380 8282 3284 8312
rect 2380 8762 3284 8792
rect 2380 9242 3284 9272
rect 2380 9722 3284 9752
rect 2380 10202 3284 10232
rect 2380 10682 3284 10712
rect 2380 11162 3284 11192
rect 2380 11642 3284 11672
rect 2380 12122 3284 12152
rect 2380 2042 2410 12152
<< m2 >>
rect 2308 1941 2390 1979
rect 2390 602 3284 640
rect 2390 1082 3284 1120
rect 2390 1562 3284 1600
rect 2390 602 2428 1979
use SUNTR_RPPO8 xa1 ../SUN_TR_SKY130NM
transform 1 0 222 0 1 222
box 222 222 2854 2340
use SUNTR_RPPO8 xa2 ../SUN_TR_SKY130NM
transform 1 0 222 0 1 2560
box 222 2560 2854 4678
use CAP_LPF xb1 
transform -1 0 20054 0 1 222
box 20054 222 36894 702
use CAP_LPF xb2_0 
transform -1 0 20054 0 1 702
box 20054 702 36894 1182
use CAP_LPF xb2_1 
transform -1 0 20054 0 1 1182
box 20054 1182 36894 1662
use CAP_LPF xb3_0 
transform -1 0 20054 0 1 1662
box 20054 1662 36894 2142
use CAP_LPF xb3_1 
transform -1 0 20054 0 1 2142
box 20054 2142 36894 2622
use CAP_LPF xb3_10 
transform -1 0 20054 0 1 2622
box 20054 2622 36894 3102
use CAP_LPF xb3_11 
transform -1 0 20054 0 1 3102
box 20054 3102 36894 3582
use CAP_LPF xb3_12 
transform -1 0 20054 0 1 3582
box 20054 3582 36894 4062
use CAP_LPF xb3_13 
transform -1 0 20054 0 1 4062
box 20054 4062 36894 4542
use CAP_LPF xb3_14 
transform -1 0 20054 0 1 4542
box 20054 4542 36894 5022
use CAP_LPF xb3_15 
transform -1 0 20054 0 1 5022
box 20054 5022 36894 5502
use CAP_LPF xb3_16 
transform -1 0 20054 0 1 5502
box 20054 5502 36894 5982
use CAP_LPF xb3_17 
transform -1 0 20054 0 1 5982
box 20054 5982 36894 6462
use CAP_LPF xb3_18 
transform -1 0 20054 0 1 6462
box 20054 6462 36894 6942
use CAP_LPF xb3_19 
transform -1 0 20054 0 1 6942
box 20054 6942 36894 7422
use CAP_LPF xb3_2 
transform -1 0 20054 0 1 7422
box 20054 7422 36894 7902
use CAP_LPF xb3_20 
transform -1 0 20054 0 1 7902
box 20054 7902 36894 8382
use CAP_LPF xb3_21 
transform -1 0 20054 0 1 8382
box 20054 8382 36894 8862
use CAP_LPF xb3_3 
transform -1 0 20054 0 1 8862
box 20054 8862 36894 9342
use CAP_LPF xb3_4 
transform -1 0 20054 0 1 9342
box 20054 9342 36894 9822
use CAP_LPF xb3_5 
transform -1 0 20054 0 1 9822
box 20054 9822 36894 10302
use CAP_LPF xb3_6 
transform -1 0 20054 0 1 10302
box 20054 10302 36894 10782
use CAP_LPF xb3_7 
transform -1 0 20054 0 1 10782
box 20054 10782 36894 11262
use CAP_LPF xb3_8 
transform -1 0 20054 0 1 11262
box 20054 11262 36894 11742
use CAP_LPF xb3_9 
transform -1 0 20054 0 1 11742
box 20054 11742 36894 12222
use cut_M1M4_2x1 xcut0 
transform 1 0 11564 0 1 0
box 11564 0 11664 38
use cut_M1M2_2x1 xcut1 
transform 1 0 530 0 1 1941
box 530 1941 622 1975
use cut_M1M2_2x1 xcut2 
transform 1 0 530 0 1 4279
box 530 4279 622 4313
use cut_M1M2_2x1 xcut3 
transform 1 0 2258 0 1 4279
box 2258 4279 2350 4313
use cut_M2M4_2x1 xcut4 
transform 1 0 3234 0 1 2042
box 3234 2042 3334 2080
use cut_M2M4_2x1 xcut5 
transform 1 0 3234 0 1 2522
box 3234 2522 3334 2560
use cut_M2M4_2x1 xcut6 
transform 1 0 3234 0 1 3002
box 3234 3002 3334 3040
use cut_M2M4_2x1 xcut7 
transform 1 0 3234 0 1 3482
box 3234 3482 3334 3520
use cut_M2M4_2x1 xcut8 
transform 1 0 3234 0 1 3962
box 3234 3962 3334 4000
use cut_M2M4_2x1 xcut9 
transform 1 0 3234 0 1 4442
box 3234 4442 3334 4480
use cut_M2M4_2x1 xcut10 
transform 1 0 3234 0 1 4922
box 3234 4922 3334 4960
use cut_M2M4_2x1 xcut11 
transform 1 0 3234 0 1 5402
box 3234 5402 3334 5440
use cut_M2M4_2x1 xcut12 
transform 1 0 3234 0 1 5882
box 3234 5882 3334 5920
use cut_M2M4_2x1 xcut13 
transform 1 0 3234 0 1 6362
box 3234 6362 3334 6400
use cut_M2M4_2x1 xcut14 
transform 1 0 3234 0 1 6842
box 3234 6842 3334 6880
use cut_M2M4_2x1 xcut15 
transform 1 0 3234 0 1 7322
box 3234 7322 3334 7360
use cut_M2M4_2x1 xcut16 
transform 1 0 3234 0 1 7802
box 3234 7802 3334 7840
use cut_M2M4_2x1 xcut17 
transform 1 0 3234 0 1 8282
box 3234 8282 3334 8320
use cut_M2M4_2x1 xcut18 
transform 1 0 3234 0 1 8762
box 3234 8762 3334 8800
use cut_M2M4_2x1 xcut19 
transform 1 0 3234 0 1 9242
box 3234 9242 3334 9280
use cut_M2M4_2x1 xcut20 
transform 1 0 3234 0 1 9722
box 3234 9722 3334 9760
use cut_M2M4_2x1 xcut21 
transform 1 0 3234 0 1 10202
box 3234 10202 3334 10240
use cut_M2M4_2x1 xcut22 
transform 1 0 3234 0 1 10682
box 3234 10682 3334 10720
use cut_M2M4_2x1 xcut23 
transform 1 0 3234 0 1 11162
box 3234 11162 3334 11200
use cut_M2M4_2x1 xcut24 
transform 1 0 3234 0 1 11642
box 3234 11642 3334 11680
use cut_M2M4_2x1 xcut25 
transform 1 0 3234 0 1 12122
box 3234 12122 3334 12160
use cut_M1M3_2x1 xcut26 
transform 1 0 2258 0 1 1941
box 2258 1941 2358 1979
use cut_M3M4_2x1 xcut27 
transform 1 0 3234 0 1 602
box 3234 602 3334 640
use cut_M3M4_2x1 xcut28 
transform 1 0 3234 0 1 1082
box 3234 1082 3334 1120
use cut_M3M4_2x1 xcut29 
transform 1 0 3234 0 1 1562
box 3234 1562 3334 1600
use cut_M1M4_1x2 xcut30 
transform 1 0 20126 0 1 0
box 20126 0 20164 100
use cut_M1M4_1x2 xcut31 
transform 1 0 20126 0 1 202
box 20126 202 20164 302
use cut_M1M4_1x2 xcut32 
transform 1 0 20126 0 1 682
box 20126 682 20164 782
use cut_M1M4_1x2 xcut33 
transform 1 0 20126 0 1 1162
box 20126 1162 20164 1262
use cut_M1M4_1x2 xcut34 
transform 1 0 20126 0 1 1642
box 20126 1642 20164 1742
use cut_M1M4_1x2 xcut35 
transform 1 0 20126 0 1 2122
box 20126 2122 20164 2222
use cut_M1M4_1x2 xcut36 
transform 1 0 20126 0 1 2602
box 20126 2602 20164 2702
use cut_M1M4_1x2 xcut37 
transform 1 0 20126 0 1 3082
box 20126 3082 20164 3182
use cut_M1M4_1x2 xcut38 
transform 1 0 20126 0 1 3562
box 20126 3562 20164 3662
use cut_M1M4_1x2 xcut39 
transform 1 0 20126 0 1 4042
box 20126 4042 20164 4142
use cut_M1M4_1x2 xcut40 
transform 1 0 20126 0 1 4522
box 20126 4522 20164 4622
use cut_M1M4_1x2 xcut41 
transform 1 0 20126 0 1 5002
box 20126 5002 20164 5102
use cut_M1M4_1x2 xcut42 
transform 1 0 20126 0 1 5482
box 20126 5482 20164 5582
use cut_M1M4_1x2 xcut43 
transform 1 0 20126 0 1 5962
box 20126 5962 20164 6062
use cut_M1M4_1x2 xcut44 
transform 1 0 20126 0 1 6442
box 20126 6442 20164 6542
use cut_M1M4_1x2 xcut45 
transform 1 0 20126 0 1 6922
box 20126 6922 20164 7022
use cut_M1M4_1x2 xcut46 
transform 1 0 20126 0 1 7402
box 20126 7402 20164 7502
use cut_M1M4_1x2 xcut47 
transform 1 0 20126 0 1 7882
box 20126 7882 20164 7982
use cut_M1M4_1x2 xcut48 
transform 1 0 20126 0 1 8362
box 20126 8362 20164 8462
use cut_M1M4_1x2 xcut49 
transform 1 0 20126 0 1 8842
box 20126 8842 20164 8942
use cut_M1M4_1x2 xcut50 
transform 1 0 20126 0 1 9322
box 20126 9322 20164 9422
use cut_M1M4_1x2 xcut51 
transform 1 0 20126 0 1 9802
box 20126 9802 20164 9902
use cut_M1M4_1x2 xcut52 
transform 1 0 20126 0 1 10282
box 20126 10282 20164 10382
use cut_M1M4_1x2 xcut53 
transform 1 0 20126 0 1 10762
box 20126 10762 20164 10862
use cut_M1M4_1x2 xcut54 
transform 1 0 20126 0 1 11242
box 20126 11242 20164 11342
use cut_M1M4_1x2 xcut55 
transform 1 0 20126 0 1 11722
box 20126 11722 20164 11822
<< labels >>
flabel locali s 20126 0 20276 12444 0 FreeSans 400 0 0 0 AVSS
port 2 nsew signal bidirectional
flabel locali s 2258 4279 2546 4389 0 FreeSans 400 0 0 0 VLPFZ
port 1 nsew signal bidirectional
flabel locali s 2258 1941 2546 2051 0 FreeSans 400 0 0 0 VLPF
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 20276 12444
<< end >>
