magic
tech sky130B
magscale 1 2
timestamp 1675206000
<< checkpaint >>
rect 0 0 2028 2880
<< locali >>
rect 1788 0 2028 2880
rect 0 0 2028 240
rect 0 2640 2028 2880
rect 0 0 240 2880
rect 1788 0 2028 2880
rect 816 530 984 590
rect 984 530 1044 590
rect 1020 678 1200 738
rect 1020 2378 1248 2438
rect 816 882 1020 942
rect 1020 678 1080 2438
rect 1140 618 1248 678
rect 1356 442 2028 502
rect 1356 794 2028 854
rect 0 516 276 576
rect 0 868 276 928
<< m2 >>
rect 1812 618 2028 678
rect 0 530 216 590
rect 1812 618 2028 678
rect 1000 618 1248 694
rect 1000 618 1920 694
rect 1000 618 1076 694
rect 0 530 216 590
rect 568 530 816 606
rect 108 530 568 606
rect 568 530 644 606
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xa2
transform 1 0 384 0 1 384
box 384 384 1644 736
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa3
transform 1 0 384 0 1 736
box 384 736 1644 2496
use cut_M1M3_2x1 
transform 1 0 1156 0 1 618
box 1156 618 1356 694
use cut_M1M3_2x1 
transform 1 0 724 0 1 530
box 724 530 924 606
<< labels >>
flabel locali s 1788 0 2028 2880 0 FreeSans 400 0 0 0 AVSS
port 3 nsew
flabel m2 s 1812 618 2028 678 0 FreeSans 400 0 0 0 IBPSR_1U
port 1 nsew
flabel m2 s 0 530 216 590 0 FreeSans 400 0 0 0 PWRUP_1V8_N
port 2 nsew
<< end >>
