magic
tech sky130B
timestamp 1728046668
<< locali >>
rect 0 2848 2172 2968
rect 0 120 120 2848
rect 192 2656 1980 2776
rect 192 312 312 2656
rect 600 2393 714 2423
rect 816 2349 1032 2379
rect 816 2173 930 2203
rect 900 2115 930 2173
rect 816 2085 930 2115
rect 585 457 615 1367
rect 1002 1323 1032 2349
rect 816 1293 1032 1323
rect 1002 443 1032 1293
rect 1590 1117 1806 1147
rect 1590 941 1704 971
rect 1674 883 1704 941
rect 1590 853 1704 883
rect 1776 707 1806 1117
rect 1590 677 1806 707
rect 1776 443 1806 677
rect 816 413 1032 443
rect 1590 413 1806 443
rect 1860 312 1980 2656
rect 192 192 1980 312
rect 2052 120 2172 2848
rect 0 0 2172 120
<< metal1 >>
rect 816 2437 930 2467
rect 816 2261 1704 2291
rect 1674 1235 1704 2261
rect 816 1205 1488 1235
rect 1590 1205 1704 1235
rect 1458 751 1488 1205
rect 1674 1059 1704 1205
rect 1590 1029 1704 1059
rect 1374 721 1488 751
rect 1458 619 1488 721
rect 1458 589 1590 619
rect 330 192 438 494
rect 762 192 870 443
rect 1104 0 1212 494
rect 1458 487 1488 589
rect 1374 457 1488 487
rect 1536 0 1644 443
<< metal2 >>
rect 816 2467 2118 2475
rect 816 2437 2172 2467
rect 54 2423 600 2431
rect 0 2393 600 2423
rect 816 2291 2118 2299
rect 816 2261 2172 2291
rect 54 2247 600 2255
rect 0 2217 600 2247
rect 54 1191 1288 1199
rect 0 1184 1288 1191
rect 0 1161 1374 1184
rect 1250 1146 1374 1161
rect 54 1015 1374 1023
rect 0 985 1374 1015
rect 54 487 600 495
rect 0 457 600 487
use SUNTR_NCHDLCM  xa1 ../SUN_TR_SKY130NM
timestamp 1728046668
transform 1 0 384 0 1 384
box -90 -66 630 946
use SUNTR_NCHDLCM  xa2
timestamp 1728046668
transform 1 0 384 0 1 1264
box -90 -66 630 946
use SUNTR_NCHDL  xa3 ../SUN_TR_SKY130NM
timestamp 1709161200
transform 1 0 384 0 1 2144
box -90 -66 630 242
use SUNTR_NCHDLA  xa4 ../SUN_TR_SKY130NM
timestamp 1728046668
transform 1 0 384 0 1 2320
box -90 -66 630 330
use SUNTR_PCHDLCM  xb1 ../SUN_TR_SKY130NM
timestamp 1728046668
transform -1 0 1788 0 1 384
box 0 -66 720 330
use SUNTR_PCHDLCM  xb2
timestamp 1728046668
transform -1 0 1788 0 1 648
box 0 -66 720 330
use SUNTR_PCHDL  xb3 ../SUN_TR_SKY130NM
timestamp 1709161200
transform -1 0 1788 0 1 912
box 0 -66 720 242
use SUNTR_PCHDL  xb4
timestamp 1709161200
transform -1 0 1788 0 1 1088
box 0 -66 720 242
use cut_M1M2_2x1  xcut0
timestamp 1720908000
transform 1 0 770 0 1 413
box 0 0 92 34
use cut_M1M2_2x1  xcut1
timestamp 1720908000
transform 1 0 770 0 1 192
box 0 0 92 34
use cut_M1M2_2x1  xcut2
timestamp 1720908000
transform 1 0 338 0 1 450
box 0 0 92 34
use cut_M1M2_2x1  xcut3
timestamp 1720908000
transform 1 0 338 0 1 192
box 0 0 92 34
use cut_M1M2_2x1  xcut4
timestamp 1720908000
transform 1 0 1544 0 1 413
box 0 0 92 34
use cut_M1M2_2x1  xcut5
timestamp 1720908000
transform 1 0 1544 0 1 0
box 0 0 92 34
use cut_M1M2_2x1  xcut6
timestamp 1720908000
transform 1 0 1112 0 1 450
box 0 0 92 34
use cut_M1M2_2x1  xcut7
timestamp 1720908000
transform 1 0 1112 0 1 0
box 0 0 92 34
use cut_M1M2_2x1  xcut8
timestamp 1720908000
transform 1 0 1320 0 1 457
box 0 0 92 34
use cut_M1M2_2x1  xcut9
timestamp 1720908000
transform 1 0 1536 0 1 589
box 0 0 92 34
use cut_M1M2_2x1  xcut10
timestamp 1720908000
transform 1 0 762 0 1 1205
box 0 0 92 34
use cut_M1M2_2x1  xcut11
timestamp 1720908000
transform 1 0 1320 0 1 721
box 0 0 92 34
use cut_M1M2_2x1  xcut12
timestamp 1720908000
transform 1 0 1536 0 1 1029
box 0 0 92 34
use cut_M1M2_2x1  xcut13
timestamp 1720908000
transform 1 0 762 0 1 2261
box 0 0 92 34
use cut_M1M2_2x1  xcut14
timestamp 1720908000
transform 1 0 1536 0 1 1205
box 0 0 92 34
use cut_M1M2_2x1  xcut15
timestamp 1720908000
transform 1 0 762 0 1 2437
box 0 0 92 34
use cut_M1M3_2x1  xcut16
timestamp 1720908000
transform 1 0 1328 0 1 1142
box 0 0 100 38
use cut_M1M3_2x1  xcut17
timestamp 1720908000
transform 1 0 554 0 1 2393
box 0 0 100 38
use cut_M1M3_2x1  xcut18
timestamp 1720908000
transform 1 0 554 0 1 457
box 0 0 100 38
use cut_M1M3_2x1  xcut19
timestamp 1720908000
transform 1 0 762 0 1 2261
box 0 0 100 38
use cut_M1M3_2x1  xcut20
timestamp 1720908000
transform 1 0 762 0 1 2437
box 0 0 100 38
use cut_M1M3_2x1  xcut21
timestamp 1720908000
transform 1 0 1328 0 1 985
box 0 0 100 38
use cut_M1M3_2x1  xcut22
timestamp 1720908000
transform 1 0 554 0 1 2217
box 0 0 100 38
<< labels >>
flabel locali s 1860 192 1980 2776 0 FreeSans 400 0 0 0 AVSS
port 6 nsew signal bidirectional
flabel locali s 2052 0 2172 2968 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel metal2 s 0 985 108 1015 0 FreeSans 400 0 0 0 CP_UP_N
port 2 nsew signal bidirectional
flabel metal2 s 2064 2261 2172 2291 0 FreeSans 400 0 0 0 LPF
port 3 nsew signal bidirectional
flabel metal2 s 0 2217 108 2247 0 FreeSans 400 0 0 0 CP_DOWN
port 4 nsew signal bidirectional
flabel metal2 s 0 457 108 487 0 FreeSans 400 0 0 0 VBN
port 5 nsew signal bidirectional
flabel metal2 s 2064 2437 2172 2467 0 FreeSans 400 0 0 0 LPFZ
port 7 nsew signal bidirectional
flabel metal2 s 0 1161 108 1191 0 FreeSans 400 0 0 0 PWRUP_1V8
port 8 nsew signal bidirectional
flabel metal2 s 0 2393 108 2423 0 FreeSans 400 0 0 0 KICK
port 9 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2172 2968
<< end >>
