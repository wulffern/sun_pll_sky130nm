magic
tech sky130B
magscale 1 2
timestamp 1675206000
<< checkpaint >>
rect 0 0 14136 7036
<< locali >>
rect 13512 384 13752 6432
rect 384 384 13752 624
rect 384 6192 13752 6432
rect 384 384 624 6432
rect 13512 384 13752 6432
rect 13896 0 14136 6816
rect 0 0 14136 240
rect 0 6576 14136 6816
rect 0 0 240 6816
rect 13896 0 14136 6816
rect 0 6960 14136 7020
rect 0 6960 14136 7020
<< m3 >>
rect 1516 384 1732 6048
rect 4844 384 5060 6048
rect 6556 384 6772 6048
rect 9884 384 10100 6048
rect 11596 384 11812 6048
rect 2308 0 2524 6048
rect 4052 0 4268 6048
rect 7348 0 7564 6048
rect 9092 0 9308 6048
rect 12388 0 12604 6048
rect 1162 4786 1238 7020
rect 5338 4786 5414 7020
rect 6202 4786 6278 7020
rect 10378 4786 10454 7020
rect 11242 4786 11318 7020
<< m1 >>
rect 1632 5578 1800 5638
rect 1800 2382 2808 2442
rect 1800 2382 1860 5638
rect 2748 2322 2856 2382
rect 6672 5578 6840 5638
rect 6840 2382 7848 2442
rect 6840 2382 6900 5638
rect 7788 2322 7896 2382
rect 11712 5578 11880 5638
rect 11880 2382 12888 2442
rect 11880 2382 11940 5638
rect 12828 2322 12936 2382
rect 4716 5578 4944 5638
rect 3768 2382 4716 2442
rect 4716 2382 4776 5638
rect 3720 2322 3828 2382
rect 9756 5578 9984 5638
rect 8808 2382 9756 2442
rect 9756 2382 9816 5638
rect 8760 2322 8868 2382
rect 1524 6960 1740 7020
rect 11172 0 11388 60
rect 11172 0 11388 60
rect 11052 1266 11280 1326
rect 11052 0 11280 60
rect 11052 0 11112 1326
rect 1524 6960 1740 7020
rect 1404 5930 1632 5990
rect 1404 6960 1632 7020
rect 1404 5930 1464 7020
<< m2 >>
rect 5376 1266 5756 1342
rect 5756 6006 6624 6082
rect 5756 1266 5832 6082
rect 6564 5930 6672 6006
rect 10416 1266 10796 1342
rect 10796 6006 11664 6082
rect 10796 1266 10872 6082
rect 11604 5930 11712 6006
rect 1248 1342 3236 1418
rect 3236 6006 4896 6082
rect 3236 1342 3312 6082
rect 1200 1266 1308 1342
rect 4836 5930 4944 6006
rect 6288 1342 8276 1418
rect 8276 6006 9936 6082
rect 8276 1342 8352 6082
rect 6240 1266 6348 1342
rect 9876 5930 9984 6006
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xc
transform 1 0 768 0 1 768
box 768 768 3288 6048
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xd
transform -1 0 5808 0 1 768
box 5808 768 8328 6048
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xe
transform 1 0 5808 0 1 768
box 5808 768 8328 6048
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xf
transform -1 0 10848 0 1 768
box 10848 768 13368 6048
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFRNQNX1_CV xg
transform 1 0 10848 0 1 768
box 10848 768 13368 6048
use cut_M1M4_2x1 
transform 1 0 1524 0 1 384
box 1524 384 1724 460
use cut_M1M4_2x1 
transform 1 0 4852 0 1 384
box 4852 384 5052 460
use cut_M1M4_2x1 
transform 1 0 6564 0 1 384
box 6564 384 6764 460
use cut_M1M4_2x1 
transform 1 0 9892 0 1 384
box 9892 384 10092 460
use cut_M1M4_2x1 
transform 1 0 11604 0 1 384
box 11604 384 11804 460
use cut_M1M4_2x1 
transform 1 0 2316 0 1 0
box 2316 0 2516 76
use cut_M1M4_2x1 
transform 1 0 4060 0 1 0
box 4060 0 4260 76
use cut_M1M4_2x1 
transform 1 0 7356 0 1 0
box 7356 0 7556 76
use cut_M1M4_2x1 
transform 1 0 9100 0 1 0
box 9100 0 9300 76
use cut_M1M4_2x1 
transform 1 0 12396 0 1 0
box 12396 0 12596 76
use cut_M2M4_2x1 
transform 1 0 1100 0 1 4786
box 1100 4786 1300 4862
use cut_M1M4_2x1 
transform 1 0 1100 0 1 6960
box 1100 6960 1300 7036
use cut_M2M4_2x1 
transform 1 0 5276 0 1 4786
box 5276 4786 5476 4862
use cut_M1M4_2x1 
transform 1 0 5276 0 1 6960
box 5276 6960 5476 7036
use cut_M2M4_2x1 
transform 1 0 6140 0 1 4786
box 6140 4786 6340 4862
use cut_M1M4_2x1 
transform 1 0 6140 0 1 6960
box 6140 6960 6340 7036
use cut_M2M4_2x1 
transform 1 0 10316 0 1 4786
box 10316 4786 10516 4862
use cut_M1M4_2x1 
transform 1 0 10316 0 1 6960
box 10316 6960 10516 7036
use cut_M2M4_2x1 
transform 1 0 11180 0 1 4786
box 11180 4786 11380 4862
use cut_M1M4_2x1 
transform 1 0 11180 0 1 6960
box 11180 6960 11380 7036
use cut_M1M2_2x1 
transform 1 0 2748 0 1 2322
box 2748 2322 2932 2390
use cut_M1M2_2x1 
transform 1 0 7788 0 1 2322
box 7788 2322 7972 2390
use cut_M1M2_2x1 
transform 1 0 12828 0 1 2322
box 12828 2322 13012 2390
use cut_M1M2_2x1 
transform 1 0 3644 0 1 2322
box 3644 2322 3828 2390
use cut_M1M2_2x1 
transform 1 0 8684 0 1 2322
box 8684 2322 8868 2390
use cut_M1M3_2x1 
transform 1 0 5268 0 1 1266
box 5268 1266 5468 1342
use cut_M1M3_2x1 
transform 1 0 6564 0 1 5930
box 6564 5930 6764 6006
use cut_M1M3_2x1 
transform 1 0 10308 0 1 1266
box 10308 1266 10508 1342
use cut_M1M3_2x1 
transform 1 0 11604 0 1 5930
box 11604 5930 11804 6006
use cut_M1M3_2x1 
transform 1 0 1092 0 1 1266
box 1092 1266 1292 1342
use cut_M1M3_2x1 
transform 1 0 4836 0 1 5930
box 4836 5930 5036 6006
use cut_M1M3_2x1 
transform 1 0 6132 0 1 1266
box 6132 1266 6332 1342
use cut_M1M3_2x1 
transform 1 0 9876 0 1 5930
box 9876 5930 10076 6006
use cut_M1M2_2x1 
transform 1 0 11204 0 1 1266
box 11204 1266 11388 1334
use cut_M1M2_2x1 
transform 1 0 1556 0 1 5930
box 1556 5930 1740 5998
<< labels >>
flabel locali s 13512 384 13752 6432 0 FreeSans 400 0 0 0 AVSS
port 5 nsew
flabel locali s 13896 0 14136 6816 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel locali s 0 6960 14136 7020 0 FreeSans 400 0 0 0 PWRUP_1V8
port 4 nsew
flabel m1 s 1524 6960 1740 7020 0 FreeSans 400 0 0 0 CK_FB
port 2 nsew
flabel m1 s 11172 0 11388 60 0 FreeSans 400 0 0 0 CK
port 3 nsew
<< end >>
