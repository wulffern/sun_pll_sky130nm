* NGSPICE file created from SUN_PLL.ext - technology: sky130B

.subckt SUNTR_NCHDL D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
C0 G B 0.412f
C1 a_324_n18# B 0.422f
C2 a_324_334# B 0.422f
.ends

.subckt SUNTR_NCHDLCM M8/a_324_334# M0/a_324_n18# D G B S
XM0 M1/S G S B M0/a_324_n18# G SUNTR_NCHDL
XM1 M2/S G M1/S B G G SUNTR_NCHDL
XM2 M3/S G M2/S B G G SUNTR_NCHDL
XM4 M5/S G M4/S B G G SUNTR_NCHDL
XM3 M4/S G M3/S B G G SUNTR_NCHDL
XM5 M6/S G M5/S B G G SUNTR_NCHDL
XM6 M7/S G M6/S B G G SUNTR_NCHDL
XM7 M8/S G M7/S B G G SUNTR_NCHDL
XM8 D G M8/S B G M8/a_324_334# SUNTR_NCHDL
C0 M8/a_324_334# B 0.422f
C1 G B 3.41f
C2 M0/a_324_n18# B 0.422f
.ends

.subckt SUN_PLL_BIAS IBPSR_1U PWRUP_1V8_N AVSS
Xxa2 IBPSR_1U PWRUP_1V8_N AVSS AVSS xa2/a_324_n18# xa2/a_324_334# SUNTR_NCHDL
Xxa3 xa3/M8/a_324_334# xa2/a_324_334# IBPSR_1U IBPSR_1U AVSS AVSS SUNTR_NCHDLCM
C0 PWRUP_1V8_N AVSS 0.884f
C1 xa3/M8/a_324_334# AVSS 0.462f
C2 IBPSR_1U AVSS 4.33f
C3 xa2/a_324_334# AVSS 0.361f
C4 xa2/a_324_n18# AVSS 0.468f
.ends

.subckt CAP_LPF A B VSUBS
R0 A m3_33320_120# sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
R1 m3_280_280# B sky130_fd_pr__res_generic_m3 w=0.4 l=0.4
C0 A B 0.232p
C1 m3_33320_120# B 0.185f
C2 m3_280_280# A 0.111f
C3 B VSUBS 48.1f
C4 A VSUBS 48.1f
.ends

.subckt SUNTR_RES8 N P a_3816_n110# a_360_n110# VSUBS
X0 a_2088_n110# a_1656_2090# VSUBS sky130_fd_pr__res_high_po w=0.72 l=8.8
X1 a_2952_n110# a_2520_2090# VSUBS sky130_fd_pr__res_high_po w=0.72 l=8.8
X2 a_2952_n110# P VSUBS sky130_fd_pr__res_high_po w=0.72 l=8.8
X3 a_360_n110# N VSUBS sky130_fd_pr__res_high_po w=0.72 l=8.8
X4 a_1224_n110# a_792_2090# VSUBS sky130_fd_pr__res_high_po w=0.72 l=8.8
X5 a_2088_n110# a_2520_2090# VSUBS sky130_fd_pr__res_high_po w=0.72 l=8.8
X6 a_360_n110# a_792_2090# VSUBS sky130_fd_pr__res_high_po w=0.72 l=8.8
X7 a_1224_n110# a_1656_2090# VSUBS sky130_fd_pr__res_high_po w=0.72 l=8.8
C0 a_2520_2090# P 0.107f
C1 a_792_2090# N 0.107f
C2 a_1656_2090# a_2520_2090# 0.107f
C3 a_792_2090# a_1656_2090# 0.107f
C4 P VSUBS 0.864f
C5 N VSUBS 0.864f
C6 a_3816_n110# VSUBS 2.55f
C7 a_2952_n110# VSUBS 0.893f
C8 a_2520_2090# VSUBS 1.1f
C9 a_2088_n110# VSUBS 0.807f
C10 a_1656_2090# VSUBS 1.1f
C11 a_1224_n110# VSUBS 0.807f
C12 a_792_2090# VSUBS 1.1f
C13 a_360_n110# VSUBS 0.893f
C14 a_n72_n110# VSUBS 2.55f $ **FLOATING
.ends

.subckt SUNTR_RPPO8 P N B XA1/a_360_n110# XA1/a_3816_n110#
XXA1 N P XA1/a_3816_n110# XA1/a_360_n110# B SUNTR_RES8
C0 P B 0.823f
C1 N B 0.823f
C2 XA1/a_3816_n110# B 2.58f
C3 XA1/a_2952_n110# B 0.936f $ **FLOATING
C4 XA1/a_2520_2090# B 1.13f $ **FLOATING
C5 XA1/a_2088_n110# B 0.838f $ **FLOATING
C6 XA1/a_1656_2090# B 1.13f $ **FLOATING
C7 XA1/a_1224_n110# B 0.838f $ **FLOATING
C8 XA1/a_792_2090# B 1.13f $ **FLOATING
C9 XA1/a_360_n110# B 0.936f
C10 XA1/a_n72_n110# B 2.58f $ **FLOATING
.ends

.subckt SUN_PLL_LPF VLPFZ VLPF AVSS
Xxb1 VLPF AVSS AVSS CAP_LPF
Xxa1 VLPF xa2/N AVSS xa1/XA1/a_360_n110# xa1/XA1/a_3816_n110# SUNTR_RPPO8
Xxa2 VLPFZ xa2/N AVSS xa2/XA1/a_360_n110# xa2/XA1/a_3816_n110# SUNTR_RPPO8
Xxb3_0 VLPFZ AVSS AVSS CAP_LPF
Xxb3_1 VLPFZ AVSS AVSS CAP_LPF
Xxb3_20 VLPFZ AVSS AVSS CAP_LPF
Xxb3_2 VLPFZ AVSS AVSS CAP_LPF
Xxb3_3 VLPFZ AVSS AVSS CAP_LPF
Xxb3_21 VLPFZ AVSS AVSS CAP_LPF
Xxb3_10 VLPFZ AVSS AVSS CAP_LPF
Xxb3_4 VLPFZ AVSS AVSS CAP_LPF
Xxb3_11 VLPFZ AVSS AVSS CAP_LPF
Xxb3_5 VLPFZ AVSS AVSS CAP_LPF
Xxb3_12 VLPFZ AVSS AVSS CAP_LPF
Xxb3_6 VLPFZ AVSS AVSS CAP_LPF
Xxb3_13 VLPFZ AVSS AVSS CAP_LPF
Xxb3_8 VLPFZ AVSS AVSS CAP_LPF
Xxb3_7 VLPFZ AVSS AVSS CAP_LPF
Xxb3_14 VLPFZ AVSS AVSS CAP_LPF
Xxb3_9 VLPFZ AVSS AVSS CAP_LPF
Xxb3_15 VLPFZ AVSS AVSS CAP_LPF
Xxb3_16 VLPFZ AVSS AVSS CAP_LPF
Xxb3_18 VLPFZ AVSS AVSS CAP_LPF
Xxb3_17 VLPFZ AVSS AVSS CAP_LPF
Xxb3_19 VLPFZ AVSS AVSS CAP_LPF
Xxb2_0 VLPF AVSS AVSS CAP_LPF
Xxb2_1 VLPF AVSS AVSS CAP_LPF
C0 VLPF VLPFZ 0.133f
C1 xa2/N xa2/XA1/a_360_n110# 0.207f
C2 xa2/XA1/a_3816_n110# VLPFZ 0.367f
C3 VLPF xa1/XA1/a_3816_n110# 0.187f
C4 VLPFZ AVSS 2.04p
C5 xa2/XA1/a_3816_n110# AVSS 2.57f
C6 xa2/XA1/a_2952_n110# AVSS 0.893f $ **FLOATING
C7 xa2/XA1/a_2520_2090# AVSS 1.1f $ **FLOATING
C8 xa2/XA1/a_2088_n110# AVSS 0.807f $ **FLOATING
C9 xa2/XA1/a_1656_2090# AVSS 1.1f $ **FLOATING
C10 xa2/XA1/a_1224_n110# AVSS 0.807f $ **FLOATING
C11 xa2/XA1/a_792_2090# AVSS 1.1f $ **FLOATING
C12 xa2/XA1/a_360_n110# AVSS 0.893f
C13 xa2/XA1/a_n72_n110# AVSS 2.56f $ **FLOATING
C14 xa2/N AVSS 3.71f
C15 xa1/XA1/a_3816_n110# AVSS 2.57f
C16 xa1/XA1/a_2952_n110# AVSS 0.893f $ **FLOATING
C17 xa1/XA1/a_2520_2090# AVSS 1.1f $ **FLOATING
C18 xa1/XA1/a_2088_n110# AVSS 0.807f $ **FLOATING
C19 xa1/XA1/a_1656_2090# AVSS 1.1f $ **FLOATING
C20 xa1/XA1/a_1224_n110# AVSS 0.807f $ **FLOATING
C21 xa1/XA1/a_792_2090# AVSS 1.1f $ **FLOATING
C22 xa1/XA1/a_360_n110# AVSS 0.893f
C23 xa1/XA1/a_n72_n110# AVSS 2.56f $ **FLOATING
C24 VLPF AVSS 0.284p
.ends

.subckt SUNTR_PCHDL D G S B a_216_n18# a_216_334# VSUBS
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
C0 B G 0.339f
C1 a_216_n18# B 0.331f
C2 a_216_334# B 0.331f
C3 B VSUBS 2.81f
.ends

.subckt SUNTR_IVX1_CV AVDD AVSS MP0/B Y MP0/a_216_n18# MP0/a_216_334# A MN0/a_324_n18#
+ VSUBS MN0/a_324_334#
XMP0 Y A AVDD MP0/B MP0/a_216_n18# MP0/a_216_334# VSUBS SUNTR_PCHDL
XMN0 Y A AVSS VSUBS MN0/a_324_n18# MN0/a_324_334# SUNTR_NCHDL
C0 MP0/B A 0.109f
C1 AVDD VSUBS 0.245f
C2 AVSS VSUBS 0.356f
C3 A VSUBS 0.628f
C4 Y VSUBS 0.264f
C5 MN0/a_324_n18# VSUBS 0.422f
C6 MN0/a_324_334# VSUBS 0.422f
C7 MP0/B VSUBS 2.81f
.ends

.subckt SUNTR_TAPCELLB_CV AVDD MN1/a_324_n18# MN1/a_324_334# MP1/a_216_334# MP1/a_216_n18#
+ AVSS
XMP1 AVDD AVDD AVDD AVDD MP1/a_216_n18# MP1/a_216_334# AVSS SUNTR_PCHDL
XMN1 AVSS AVSS AVSS AVSS MN1/a_324_n18# MN1/a_324_334# SUNTR_NCHDL
C0 AVDD AVSS 0.105f
C1 AVSS 0 1.04f
C2 MN1/a_324_n18# 0 0.422f
C3 MN1/a_324_334# 0 0.422f
C4 AVDD 0 3.14f
.ends

.subckt SUNTR_DFTSPCX1_CV CK Q AVDD AVSS MN1/a_324_334# MP2/B D MP2/G MP1/a_216_n18#
+ MN0/a_324_n18# MP2/a_216_334# VSUBS
XMP0 MP2/G CK MP1/D MP2/B MP1/a_216_334# MP2/a_216_n18# VSUBS SUNTR_PCHDL
XMP1 MP1/D D AVDD MP2/B MP1/a_216_n18# MP1/a_216_334# VSUBS SUNTR_PCHDL
XMP2 Q MP2/G AVDD MP2/B MP2/a_216_n18# MP2/a_216_334# VSUBS SUNTR_PCHDL
XMN0 MP2/G D AVSS VSUBS MN0/a_324_n18# MN2/a_324_n18# SUNTR_NCHDL
XMN1 AVSS MP2/G MN2/D VSUBS MN2/a_324_334# MN1/a_324_334# SUNTR_NCHDL
XMN2 MN2/D CK Q VSUBS MN2/a_324_n18# MN2/a_324_334# SUNTR_NCHDL
C0 MP2/B MP2/a_216_n18# -0.311f
C1 MP1/a_216_334# MP2/B -0.311f
C2 MP2/G AVDD 0.102f
C3 MP2/G Q 0.241f
C4 MP2/G CK 0.173f
C5 MP2/B AVDD 0.211f
C6 MP2/B CK 0.111f
C7 AVSS AVDD 0.132f
C8 MP2/B D 0.11f
C9 MP2/B MP2/G 0.211f
C10 AVDD VSUBS 0.343f
C11 AVSS VSUBS 0.602f
C12 Q VSUBS 0.242f
C13 CK VSUBS 0.477f
C14 MN2/a_324_n18# VSUBS 0.35f
C15 MN2/a_324_334# VSUBS 0.35f
C16 MN1/a_324_334# VSUBS 0.422f
C17 D VSUBS 0.551f
C18 MP2/G VSUBS 1.15f
C19 MN0/a_324_n18# VSUBS 0.422f
C20 MP2/B VSUBS 5.96f
.ends

.subckt SUNTR_NRX1_CV B AVDD AVSS MN1/a_324_334# MP1/B A MP0/a_216_n18# Y MP1/a_216_334#
+ MN0/a_324_n18# VSUBS
XMP0 MP1/S A AVDD MP1/B MP0/a_216_n18# MP1/a_216_n18# VSUBS SUNTR_PCHDL
XMP1 Y B MP1/S MP1/B MP1/a_216_n18# MP1/a_216_334# VSUBS SUNTR_PCHDL
XMN0 Y A AVSS VSUBS MN0/a_324_n18# MN1/a_324_n18# SUNTR_NCHDL
XMN1 AVSS B Y VSUBS MN1/a_324_n18# MN1/a_324_334# SUNTR_NCHDL
C0 MP1/a_216_n18# MP1/B -0.311f
C1 AVDD MP1/B 0.136f
C2 Y AVSS 0.122f
C3 MP1/B B 0.11f
C4 MP1/B A 0.11f
C5 AVSS VSUBS 0.54f
C6 Y VSUBS 0.306f
C7 B VSUBS 0.561f
C8 MN1/a_324_n18# VSUBS 0.353f
C9 MN1/a_324_334# VSUBS 0.422f
C10 A VSUBS 0.562f
C11 MN0/a_324_n18# VSUBS 0.422f
C12 MP1/B VSUBS 4.38f
C13 AVDD VSUBS 0.269f
.ends

.subckt SUN_PLL_PFD CP_UP_N CK_REF CP_DOWN CK_FB AVDD xa5/D AVSS
Xxa2a AVDD AVSS AVDD CP_UP_N xa2/MP0/a_216_334# xa3/MP0/a_216_n18# xa2/Y xa2/MN0/a_324_334#
+ AVSS xa3/MN0/a_324_n18# SUNTR_IVX1_CV
Xxa0 AVDD xa0/MN1/a_324_n18# xa1/MN0/a_324_n18# xa1/MP1/a_216_n18# xa0/MP1/a_216_n18#
+ AVSS SUNTR_TAPCELLB_CV
Xxa1 CK_REF xa3/A AVDD AVSS xa2/MN0/a_324_n18# AVDD xa5/D xa1/MP2/G xa1/MP1/a_216_n18#
+ xa1/MN0/a_324_n18# xa2/MP0/a_216_n18# AVSS SUNTR_DFTSPCX1_CV
Xxa2 AVDD AVSS AVDD xa2/Y xa2/MP0/a_216_n18# xa2/MP0/a_216_334# xa3/A xa2/MN0/a_324_n18#
+ AVSS xa2/MN0/a_324_334# SUNTR_IVX1_CV
Xxa3 xa6/A AVDD AVSS xa5/MN0/a_324_n18# AVDD xa3/A xa3/MP0/a_216_n18# xa5/D xa5/MP1/a_216_n18#
+ xa3/MN0/a_324_n18# AVSS SUNTR_NRX1_CV
Xxa5 CK_FB xa6/A AVDD AVSS xa6/MN0/a_324_n18# AVDD xa5/D xa5/MP2/G xa5/MP1/a_216_n18#
+ xa5/MN0/a_324_n18# xa6/MP0/a_216_n18# AVSS SUNTR_DFTSPCX1_CV
Xxa6 AVDD AVSS AVDD CP_DOWN xa6/MP0/a_216_n18# xa6/MP0/a_216_334# xa6/A xa6/MN0/a_324_n18#
+ AVSS xa6/MN0/a_324_334# SUNTR_IVX1_CV
C0 AVSS xa3/A 0.157f
C1 AVDD xa2/MP0/a_216_n18# -0.311f
C2 AVDD xa5/D 0.14f
C3 xa5/D xa6/A 0.344f
C4 xa2/Y xa3/A 0.342f
C5 AVSS CP_DOWN 0.482f
C6 AVDD xa3/MP0/a_216_n18# -0.313f
C7 AVDD xa6/MP0/a_216_n18# -0.312f
C8 AVDD xa1/MP1/a_216_n18# -0.311f
C9 AVDD AVSS 5.16f
C10 xa6/A xa5/MP2/G 0.195f
C11 AVSS xa6/A 0.314f
C12 xa2/Y AVSS 0.201f
C13 CP_UP_N AVSS 0.451f
C14 AVDD CP_DOWN 0.539f
C15 AVDD xa6/A 0.113f
C16 CP_UP_N AVDD 0.697f
C17 xa1/MP2/G xa5/D 0.179f
C18 AVSS CK_REF 0.179f
C19 xa3/A xa1/MP2/G 0.171f
C20 AVDD xa5/MP1/a_216_n18# -0.311f
C21 AVDD xa2/MP0/a_216_334# -0.311f
C22 AVSS xa5/D 0.515f
C23 AVSS CK_FB 0.178f
C24 CP_DOWN 0 0.516f
C25 xa6/MN0/a_324_n18# 0 0.36f
C26 xa6/MN0/a_324_334# 0 0.422f
C27 CK_FB 0 0.773f
C28 xa5/MN2/a_324_n18# 0 0.355f
C29 xa5/MN2/a_324_334# 0 0.355f
C30 xa5/MP2/G 0 1.03f
C31 xa5/MN0/a_324_n18# 0 0.36f
C32 xa6/A 0 1.62f
C33 xa3/MN1/a_324_n18# 0 0.355f
C34 xa3/MN0/a_324_n18# 0 0.36f
C35 xa3/A 0 1.5f
C36 xa2/MN0/a_324_n18# 0 0.36f
C37 xa2/MN0/a_324_334# 0 0.36f
C38 CK_REF 0 0.768f
C39 xa1/MN2/a_324_n18# 0 0.355f
C40 xa1/MN2/a_324_334# 0 0.355f
C41 xa5/D 0 1.97f
C42 xa1/MP2/G 0 1.03f
C43 xa1/MN0/a_324_n18# 0 0.36f
C44 AVSS 0 1.63f
C45 xa0/MN1/a_324_n18# 0 0.422f
C46 AVDD 0 29.2f
C47 xa2/Y 0 0.716f
C48 CP_UP_N 0 0.39f
.ends

.subckt SUNTR_PCHDLCM M7/a_216_334# D G M0/a_216_n18# B VSUBS S
XM0 M7/S G S B M0/a_216_n18# G VSUBS SUNTR_PCHDL
XM7 D G M7/S B G M7/a_216_334# VSUBS SUNTR_PCHDL
C0 B G -0.658f
C1 G VSUBS 0.104f
C2 B VSUBS 3.6f
.ends

.subckt SUNTR_NCHDLA G D M0/a_324_n18# B S
XM0 D G S B M0/a_324_n18# G SUNTR_NCHDL
XM1 S G D B G M1/a_324_334# SUNTR_NCHDL
C0 M1/a_324_334# B 0.422f
C1 S B 0.285f
C2 G B 0.776f
C3 M0/a_324_n18# B 0.422f
.ends

.subckt SUN_PLL_CP AVDD CP_UP_N LPF CP_DOWN VBN LPFZ PWRUP_1V8 KICK AVSS
Xxb1 xb2/M0/a_216_n18# xb2/G xb2/G xb1/M0/a_216_n18# AVDD AVSS AVDD SUNTR_PCHDLCM
Xxb2 xb3/a_216_n18# xb3/S xb2/G xb2/M0/a_216_n18# AVDD AVSS AVDD SUNTR_PCHDLCM
Xxa1 xa2/M0/a_324_n18# xa1/M0/a_324_n18# xb2/G VBN AVSS AVSS SUNTR_NCHDLCM
Xxa2 xa3/a_324_n18# xa2/M0/a_324_n18# xa3/S VBN AVSS AVSS SUNTR_NCHDLCM
Xxb3 LPF CP_UP_N xb3/S AVDD xb3/a_216_n18# xb4/a_216_n18# AVSS SUNTR_PCHDL
Xxa3 LPF CP_DOWN xa3/S AVSS xa3/a_324_n18# xa3/a_324_334# SUNTR_NCHDL
Xxb4 LPF PWRUP_1V8 AVDD AVDD xb4/a_216_n18# xb4/a_216_334# AVSS SUNTR_PCHDL
Xxa4 KICK LPFZ xa3/a_324_334# AVSS AVSS SUNTR_NCHDLA
C0 KICK CP_DOWN 0.239f
C1 xb2/G PWRUP_1V8 0.249f
C2 AVDD xb4/a_216_n18# -0.302f
C3 LPFZ LPF 0.477f
C4 VBN CP_UP_N 0.139f
C5 xb3/S AVDD 0.105f
C6 VBN AVDD 0.122f
C7 CP_UP_N PWRUP_1V8 0.479f
C8 xb3/a_216_n18# AVDD -0.31f
C9 xb2/G AVDD 0.852f
C10 AVDD PWRUP_1V8 0.203f
C11 AVDD LPF 0.369f
C12 AVDD xb2/M0/a_216_n18# -0.302f
C13 AVDD CP_UP_N 0.247f
C14 PWRUP_1V8 AVSS 0.603f
C15 CP_DOWN AVSS 0.735f
C16 LPF AVSS 2.37f
C17 xa4/M1/a_324_334# AVSS 0.461f
C18 KICK AVSS 1.15f
C19 LPFZ AVSS 0.793f
C20 xa3/a_324_334# AVSS 0.358f
C21 xa3/S AVSS 0.166f
C22 xa3/a_324_n18# AVSS 0.356f
C23 xa2/M0/a_324_n18# AVSS 0.36f
C24 VBN AVSS 7.29f
C25 xa1/M0/a_324_n18# AVSS 0.494f
C26 xb2/G AVSS 0.736f
C27 AVDD AVSS 18.1f
C28 xb1/M0/a_216_n18# AVSS 0.131f
C29 CP_UP_N AVSS 0.44f
.ends

.subckt SUNTR_DCAPX1_CV A B li_2412_n44# li_n108_n44# VSUBS
R0 li_468_484# B sky130_fd_pr__res_generic_l1 w=0.44 l=0.36
R1 A li_1836_1012# sky130_fd_pr__res_generic_l1 w=0.44 l=0.36
C0 B A 1.75f
C1 B li_2412_n44# 0.111f
C2 B li_1836_1012# 0.117f
C3 li_n108_n44# A 0.108f
C4 B VSUBS 1.23f
C5 A VSUBS 1.85f
C6 li_2412_n44# VSUBS 0.968f
C7 li_n108_n44# VSUBS 0.979f
.ends

.subckt SUN_PLL_KICK KICK KICK_N PWRUP_1V8_N AVDD AVSS PWRUP_1V8
Xxa5a AVDD AVSS AVDD xa6/A xa2/MP0/a_216_334# xa5a/MP0/a_216_334# xa2/Y xa2/MN0/a_324_334#
+ AVSS xa5a/MN0/a_324_334# SUNTR_IVX1_CV
Xxa1a AVDD xa1a/MN1/a_324_n18# xa1b/MN0/a_324_n18# xa1b/MP0/a_216_n18# xa1a/MP1/a_216_n18#
+ AVSS SUNTR_TAPCELLB_CV
Xxa1b AVDD AVSS AVDD PWRUP_1V8_N xa1b/MP0/a_216_n18# xa1c/MP0/a_216_n18# PWRUP_1V8
+ xa1b/MN0/a_324_n18# AVSS xa1c/MN0/a_324_n18# SUNTR_IVX1_CV
Xxa1c AVDD AVSS AVDD xa2/A xa1c/MP0/a_216_n18# xa2/MP0/a_216_n18# PWRUP_1V8_N xa1c/MN0/a_324_n18#
+ AVSS xa2/MN0/a_324_n18# SUNTR_IVX1_CV
Xxa2 AVDD AVSS AVDD xa2/Y xa2/MP0/a_216_n18# xa2/MP0/a_216_334# xa2/A xa2/MN0/a_324_n18#
+ AVSS xa2/MN0/a_324_334# SUNTR_IVX1_CV
Xxa6 AVDD AVSS AVDD xa7/A xa6/MP0/a_216_n18# xa7/MP0/a_216_n18# xa6/A xa6/MN0/a_324_n18#
+ AVSS xa7/MN0/a_324_n18# SUNTR_IVX1_CV
Xxa7 AVDD AVSS AVDD xa8/B xa7/MP0/a_216_n18# xa8/MP0/a_216_n18# xa7/A xa7/MN0/a_324_n18#
+ AVSS xa8/MN0/a_324_n18# SUNTR_IVX1_CV
Xxa8 xa8/B AVDD AVSS xa9/MN0/a_324_n18# AVDD PWRUP_1V8_N xa8/MP0/a_216_n18# KICK xa9/MP0/a_216_n18#
+ xa8/MN0/a_324_n18# AVSS SUNTR_NRX1_CV
Xxa9 AVDD AVSS AVDD KICK_N xa9/MP0/a_216_n18# xa9/MP0/a_216_334# KICK xa9/MN0/a_324_n18#
+ AVSS xa9/MN0/a_324_334# SUNTR_IVX1_CV
Xxa5capb AVSS xa6/A AVDD AVSS AVSS SUNTR_DCAPX1_CV
C0 AVDD xa7/MP0/a_216_n18# -0.311f
C1 AVDD xa2/MP0/a_216_n18# -0.311f
C2 AVSS xa2/A 0.238f
C3 AVDD PWRUP_1V8_N 0.108f
C4 AVSS KICK 0.218f
C5 AVDD AVSS 5.06f
C6 xa6/A xa2/Y 0.113f
C7 xa6/A xa7/A 0.124f
C8 AVSS KICK_N 0.114f
C9 AVDD xa1c/MP0/a_216_n18# -0.311f
C10 PWRUP_1V8_N xa6/A 0.225f
C11 AVSS xa8/B 0.151f
C12 PWRUP_1V8_N xa7/A 0.137f
C13 AVSS xa2/Y 0.253f
C14 AVSS xa6/A 0.847f
C15 AVDD xa1b/MP0/a_216_n18# -0.311f
C16 AVSS xa7/A 0.28f
C17 AVDD xa2/MP0/a_216_334# -0.311f
C18 xa8/B KICK 0.25f
C19 xa2/Y xa2/A 0.182f
C20 AVDD xa9/MP0/a_216_n18# -0.311f
C21 PWRUP_1V8_N PWRUP_1V8 0.108f
C22 AVDD xa6/A 0.367f
C23 AVDD xa8/MP0/a_216_n18# -0.311f
C24 AVSS PWRUP_1V8_N 0.879f
C25 PWRUP_1V8_N xa2/A 0.215f
C26 xa9/MN0/a_324_334# 0 0.422f
C27 KICK 0 0.897f
C28 xa8/MN1/a_324_n18# 0 0.355f
C29 xa9/MN0/a_324_n18# 0 0.36f
C30 xa8/MN0/a_324_n18# 0 0.36f
C31 xa8/B 0 0.768f
C32 xa7/MN0/a_324_n18# 0 0.36f
C33 xa7/A 0 0.716f
C34 xa6/MN0/a_324_n18# 0 0.422f
C35 xa2/MN0/a_324_n18# 0 0.36f
C36 xa2/A 0 0.703f
C37 xa1c/MN0/a_324_n18# 0 0.36f
C38 PWRUP_1V8 0 0.512f
C39 PWRUP_1V8_N 0 2.14f
C40 xa1b/MN0/a_324_n18# 0 0.36f
C41 AVSS 0 4.7f
C42 xa1a/MN1/a_324_n18# 0 0.422f
C43 AVDD 0 29.1f
C44 xa2/Y 0 0.756f
C45 xa6/A 0 2.53f
C46 xa2/MN0/a_324_334# 0 0.36f
C47 xa5a/MN0/a_324_334# 0 0.422f
.ends

.subckt SUNSAR_CAP_BSSW_CV A B VSUBS
R0 A m3_9828_132# sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
R1 m3_252_308# B sky130_fd_pr__res_generic_m3 w=0.44 l=0.36
C0 A B 64.5f
C1 m3_9828_132# B 0.17f
C2 m3_252_308# A 0.106f
C3 B VSUBS 15.7f
C4 A VSUBS 15.7f
.ends

.subckt SUNTR_PCHL D G S B a_216_492# a_216_n36# VSUBS
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.518 pd=3.12 as=0.518 ps=3.12 w=1.08 l=0.36
C0 B G 0.398f
C1 a_216_n36# B 0.426f
C2 a_216_492# B 0.427f
C3 B VSUBS 3.6f
C4 a_216_n36# VSUBS 0.106f
C5 a_216_492# VSUBS 0.106f
.ends

.subckt SUN_PLL_BUF AVDD VFB VI VO VBN AVSS
Xxd3_0 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxd3_1 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxd3_2 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxd3_3 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxd3_5 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxc3_11 VO xc3_9/G AVDD AVDD xc3_12/a_216_n36# xc3_11/a_216_n36# AVSS SUNTR_PCHL
Xxd3_4 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxc3_10 VO xc3_9/G AVDD AVDD xc3_11/a_216_n36# xc3_1/a_216_492# AVSS SUNTR_PCHL
Xxd3_6 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxc3_12 VO xc3_9/G AVDD AVDD xc3_2/a_216_n36# xc3_12/a_216_n36# AVSS SUNTR_PCHL
Xxd3_7 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxd3_8 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxc2_1 xc3_9/G xc2_3/G AVDD AVDD xc2_2/a_216_n36# xc2_1/a_216_n36# AVSS SUNTR_PCHL
Xxc2_0 xc3_9/G xc2_3/G AVDD AVDD xc2_1/a_216_n36# xc2_0/a_216_n36# AVSS SUNTR_PCHL
Xxd3_9 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxc2_2 xc3_9/G xc2_3/G AVDD AVDD xc2_3/a_216_n36# xc2_2/a_216_n36# AVSS SUNTR_PCHL
Xxd2 VO AVSS AVSS SUNSAR_CAP_BSSW_CV
Xxc2_3 xc3_9/G xc2_3/G AVDD AVDD xc3_0/a_216_n36# xc2_3/a_216_n36# AVSS SUNTR_PCHL
Xxa1 xa1/M8/a_324_334# xa1/M0/a_324_n18# xa1/D VBN AVSS AVSS SUNTR_NCHDLCM
Xxa4_0 xa4_1/M0/a_324_n18# xa4_0/M0/a_324_n18# xc3_9/G VI AVSS xa1/D SUNTR_NCHDLCM
Xxa4_1 xa4_1/M8/a_324_334# xa4_1/M0/a_324_n18# xc3_9/G VI AVSS xa1/D SUNTR_NCHDLCM
Xxa2_0 xa2_1/M0/a_324_n18# xa1/M8/a_324_334# xc2_3/G VFB AVSS xa1/D SUNTR_NCHDLCM
Xxa2_1 xa4_0/M0/a_324_n18# xa2_1/M0/a_324_n18# xc2_3/G VFB AVSS xa1/D SUNTR_NCHDLCM
Xxc3_0 VO xc3_9/G AVDD AVDD xc3_1/a_216_n36# xc3_0/a_216_n36# AVSS SUNTR_PCHL
Xxc3_1 VO xc3_9/G AVDD AVDD xc3_1/a_216_492# xc3_1/a_216_n36# AVSS SUNTR_PCHL
Xxc3_2 VO xc3_9/G AVDD AVDD xc3_3/a_216_n36# xc3_2/a_216_n36# AVSS SUNTR_PCHL
Xxc3_3 VO xc3_9/G AVDD AVDD xc3_4/a_216_n36# xc3_3/a_216_n36# AVSS SUNTR_PCHL
Xxc1_0 xc2_3/G xc2_3/G AVDD AVDD xc1_1/a_216_n36# xc1_0/a_216_n36# AVSS SUNTR_PCHL
Xxc3_4 VO xc3_9/G AVDD AVDD xc3_5/a_216_n36# xc3_4/a_216_n36# AVSS SUNTR_PCHL
Xxc1_1 xc2_3/G xc2_3/G AVDD AVDD xc1_2/a_216_n36# xc1_1/a_216_n36# AVSS SUNTR_PCHL
Xxc3_5 VO xc3_9/G AVDD AVDD xc3_6/a_216_n36# xc3_5/a_216_n36# AVSS SUNTR_PCHL
Xxc1_2 xc2_3/G xc2_3/G AVDD AVDD xc1_3/a_216_n36# xc1_2/a_216_n36# AVSS SUNTR_PCHL
Xxc3_7 VO xc3_9/G AVDD AVDD xc3_8/a_216_n36# xc3_7/a_216_n36# AVSS SUNTR_PCHL
Xxc3_6 VO xc3_9/G AVDD AVDD xc3_7/a_216_n36# xc3_6/a_216_n36# AVSS SUNTR_PCHL
Xxc1_3 xc2_3/G xc2_3/G AVDD AVDD xc2_0/a_216_n36# xc1_3/a_216_n36# AVSS SUNTR_PCHL
Xxc3_8 VO xc3_9/G AVDD AVDD xc3_9/a_216_n36# xc3_8/a_216_n36# AVSS SUNTR_PCHL
Xxc3_9 VO xc3_9/G AVDD AVDD xc3_9/a_216_492# xc3_9/a_216_n36# AVSS SUNTR_PCHL
C0 xc3_5/a_216_n36# AVDD -0.349f
C1 xc2_3/a_216_n36# AVDD -0.349f
C2 xc3_11/a_216_n36# AVDD -0.349f
C3 xc1_1/a_216_n36# AVDD -0.347f
C4 VO xc2_3/G 0.573f
C5 VO AVDD 5.72f
C6 AVDD xc2_3/G 2.56f
C7 VI VFB 0.212f
C8 VO xc3_9/G 1.26f
C9 xc3_1/a_216_n36# AVDD -0.349f
C10 xc3_9/G xc2_3/G 0.709f
C11 xc3_9/G AVDD 4.1f
C12 xc2_2/a_216_n36# AVDD -0.349f
C13 xa1/D VI 0.182f
C14 xc3_9/a_216_n36# AVDD -0.349f
C15 xa1/D VFB 0.372f
C16 xc3_8/a_216_n36# AVDD -0.349f
C17 xc3_12/a_216_n36# AVDD -0.349f
C18 xc3_3/a_216_n36# AVDD -0.349f
C19 xc1_3/a_216_n36# AVDD -0.349f
C20 xc3_2/a_216_n36# AVDD -0.349f
C21 VI AVDD 0.246f
C22 xc2_0/a_216_n36# AVDD -0.349f
C23 xc3_6/a_216_n36# AVDD -0.349f
C24 VFB AVDD 0.411f
C25 xc2_1/a_216_n36# AVDD -0.349f
C26 xc3_7/a_216_n36# AVDD -0.349f
C27 xa1/D xc2_3/G 0.238f
C28 xc3_1/a_216_492# AVDD -0.349f
C29 xa1/D AVDD 0.321f
C30 xc1_2/a_216_n36# AVDD -0.349f
C31 VBN AVDD 0.148f
C32 xc3_4/a_216_n36# AVDD -0.349f
C33 xa1/D xc3_9/G 0.141f
C34 xc3_0/a_216_n36# AVDD -0.349f
C35 xc2_3/G AVSS 1.65f
C36 AVDD AVSS 65.4f
C37 xc3_9/G AVSS 2.08f
C38 xc3_9/a_216_492# AVSS 0.11f
C39 xc1_0/a_216_n36# AVSS 0.17f
C40 xa4_0/M0/a_324_n18# AVSS 0.354f
C41 xa2_1/M0/a_324_n18# AVSS 0.353f
C42 VFB AVSS 8.32f
C43 xa1/M8/a_324_334# AVSS 0.354f
C44 xa4_1/M8/a_324_334# AVSS 0.422f
C45 xa4_1/M0/a_324_n18# AVSS 0.353f
C46 VI AVSS 7.32f
C47 xa1/D AVSS 1.44f
C48 VBN AVSS 3.86f
C49 xa1/M0/a_324_n18# AVSS 0.488f
C50 VO AVSS 0.277p
.ends

.subckt SUNTRB_PCHDL D G S B a_216_n18# a_216_334# VSUBS
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
C0 a_216_n18# B 0.331f
C1 a_216_334# B 0.331f
C2 B G 0.339f
C3 B VSUBS 2.81f
.ends

.subckt SUNTRB_NCHDL D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.616 pd=3.3 as=0.616 ps=3.3 w=1.08 l=0.18
C0 G B 0.412f
C1 a_324_n18# B 0.422f
C2 a_324_334# B 0.422f
.ends

.subckt SUNTRB_IVX1_CV BULKP AVDD AVSS A Y MP0/a_216_n18# MP0/a_216_334# MN0/a_324_n18#
+ VSUBS MN0/a_324_334#
XMP0 Y A AVDD BULKP MP0/a_216_n18# MP0/a_216_334# VSUBS SUNTRB_PCHDL
XMN0 Y A AVSS VSUBS MN0/a_324_n18# MN0/a_324_334# SUNTRB_NCHDL
C0 BULKP A 0.109f
C1 AVSS VSUBS 0.356f
C2 Y VSUBS 0.264f
C3 MN0/a_324_n18# VSUBS 0.422f
C4 MN0/a_324_334# VSUBS 0.422f
C5 AVDD VSUBS 0.245f
C6 A VSUBS 0.628f
C7 BULKP VSUBS 2.81f
.ends

.subckt SUNTRB_NDX1_CV B Y AVDD AVSS MN1/a_324_334# A BULKP MP1/a_216_334# VSUBS
XMP0 Y A AVDD BULKP MP0/a_216_n18# MP1/a_216_n18# VSUBS SUNTRB_PCHDL
XMP1 AVDD B Y BULKP MP1/a_216_n18# MP1/a_216_334# VSUBS SUNTRB_PCHDL
XMN0 MN1/S A AVSS VSUBS MN0/a_324_n18# MN1/a_324_n18# SUNTRB_NCHDL
XMN1 Y B MN1/S VSUBS MN1/a_324_n18# MN1/a_324_334# SUNTRB_NCHDL
C0 BULKP AVDD 0.175f
C1 BULKP Y 0.115f
C2 BULKP B 0.11f
C3 A BULKP 0.11f
C4 MP1/a_216_n18# BULKP -0.311f
C5 AVSS VSUBS 0.411f
C6 MN1/a_324_334# VSUBS 0.422f
C7 AVDD VSUBS 0.345f
C8 MN0/a_324_n18# VSUBS 0.422f
C9 MN1/a_324_n18# VSUBS 0.352f
C10 Y VSUBS 0.299f
C11 B VSUBS 0.561f
C12 BULKP VSUBS 4.38f
C13 A VSUBS 0.562f
.ends

.subckt SUNTRB_TAPCELLBAVSS_CV MN1/a_324_n18# MP1/B MP1/a_216_n18# AVSS
XMP1 MP1/S MP1/S MP1/S MP1/B MP1/a_216_n18# MP1/a_216_334# AVSS SUNTRB_PCHDL
XMN1 AVSS AVSS AVSS AVSS MN1/a_324_n18# MN1/a_324_334# SUNTRB_NCHDL
C0 AVSS 0 1.07f
C1 MN1/a_324_n18# 0 0.422f
C2 MN1/a_324_334# 0 0.422f
C3 MP1/S 0 0.177f
C4 MP1/B 0 2.81f
.ends

.subckt SUN_PLL_LSCORE A AVDD AVSS xb2_1/a_324_334# xc2b/a_216_334# YN xc2b/B AN Y
+ VSUBS
Xxc2a xc2b/S Y AVDD xc2b/B xc2a/a_216_n18# xc2b/a_216_n18# VSUBS SUNTR_PCHDL
Xxc2b YN Y xc2b/S xc2b/B xc2b/a_216_n18# xc2b/a_216_334# VSUBS SUNTR_PCHDL
Xxc1a xc1b/S YN AVDD xc2b/B xc1a/a_216_n18# xc1b/a_216_n18# VSUBS SUNTR_PCHDL
Xxc1b Y YN xc1b/S xc2b/B xc1b/a_216_n18# xc2a/a_216_n18# VSUBS SUNTR_PCHDL
Xxb1_0 Y AN AVSS VSUBS xb1_0/a_324_n18# xb1_1/a_324_n18# SUNTR_NCHDL
Xxb1_1 Y AN AVSS VSUBS xb1_1/a_324_n18# xb2_0/a_324_n18# SUNTR_NCHDL
Xxb2_0 YN A AVSS VSUBS xb2_0/a_324_n18# xb2_1/a_324_n18# SUNTR_NCHDL
Xxb2_1 YN A AVSS VSUBS xb2_1/a_324_n18# xb2_1/a_324_334# SUNTR_NCHDL
C0 Y AVSS 0.224f
C1 xc2a/a_216_n18# xc2b/B -0.311f
C2 xc2b/B Y 0.334f
C3 YN AVSS 0.161f
C4 YN Y 0.347f
C5 AVSS AVDD 0.185f
C6 Y AVDD 0.253f
C7 xc1b/a_216_n18# xc2b/B -0.311f
C8 YN xc2b/B 0.414f
C9 xc2b/a_216_n18# xc2b/B -0.311f
C10 xc2b/B AVDD 0.222f
C11 AVDD VSUBS 0.362f
C12 xb2_1/a_324_n18# VSUBS 0.352f
C13 xb2_1/a_324_334# VSUBS 0.422f
C14 A VSUBS 0.874f
C15 xb2_0/a_324_n18# VSUBS 0.353f
C16 xb1_1/a_324_n18# VSUBS 0.352f
C17 AVSS VSUBS 0.742f
C18 AN VSUBS 0.874f
C19 Y VSUBS 0.435f
C20 xb1_0/a_324_n18# VSUBS 0.422f
C21 xc2b/B VSUBS 7.54f
C22 YN VSUBS 0.421f
.ends

.subckt SUN_PLL_ROSC AVDD CK VDD_ROSC PWRUP_1V8 AVSS
Xxb2_3 AVDD VDD_ROSC AVSS xb2_3/A xb2_4/A xb2_3/MP0/a_216_n18# xb2_4/MP0/a_216_n18#
+ xb2_3/MN0/a_324_n18# AVSS xb2_4/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_2 AVDD VDD_ROSC AVSS xb2_2/A xb2_3/A xb2_2/MP0/a_216_n18# xb2_3/MP0/a_216_n18#
+ xb2_2/MN0/a_324_n18# AVSS xb2_3/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_4 AVDD VDD_ROSC AVSS xb2_4/A xb2_5/A xb2_4/MP0/a_216_n18# xb2_5/MP0/a_216_n18#
+ xb2_4/MN0/a_324_n18# AVSS xb2_5/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_5 AVDD VDD_ROSC AVSS xb2_5/A xa3/A xb2_5/MP0/a_216_n18# xb2_6/MP0/a_216_n18#
+ xb2_5/MN0/a_324_n18# AVSS xb2_6/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_6 AVDD VDD_ROSC AVSS xa3/A xa3/AN xb2_6/MP0/a_216_n18# xb2_7/MP0/a_216_n18# xb2_6/MN0/a_324_n18#
+ AVSS xb2_7/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_7 AVDD VDD_ROSC AVSS xa3/AN xb1/B xb2_7/MP0/a_216_n18# xb3/MP1/a_216_n18# xb2_7/MN0/a_324_n18#
+ AVSS xb3/MN1/a_324_n18# SUNTRB_IVX1_CV
Xxb1 xb1/B xb1/Y VDD_ROSC AVSS xb1/MN1/a_324_334# PWRUP_1V8 AVDD xb1/MP1/a_216_334#
+ AVSS SUNTRB_NDX1_CV
Xxb3 xb3/MN1/a_324_n18# AVDD xb3/MP1/a_216_n18# AVSS SUNTRB_TAPCELLBAVSS_CV
Xxa3 xa3/A AVDD AVSS xa4/MN0/a_324_n18# xa4/MP0/a_216_n18# xa5/A AVDD xa3/AN xa4/A
+ AVSS SUN_PLL_LSCORE
Xxa4 AVDD AVSS AVDD xa4/Y xa4/MP0/a_216_n18# xa5/MP0/a_216_n18# xa4/A xa4/MN0/a_324_n18#
+ AVSS xa5/MN0/a_324_n18# SUNTR_IVX1_CV
Xxa5 AVDD AVSS AVDD CK xa5/MP0/a_216_n18# xa6/MP1/a_216_n18# xa5/A xa5/MN0/a_324_n18#
+ AVSS xa6/MN1/a_324_n18# SUNTR_IVX1_CV
Xxa6 AVDD xa6/MN1/a_324_n18# xa6/MN1/a_324_334# xa6/MP1/a_216_334# xa6/MP1/a_216_n18#
+ AVSS SUNTR_TAPCELLB_CV
Xxb2_0 AVDD VDD_ROSC AVSS xb1/Y xb2_1/A xb1/MP1/a_216_334# xb2_1/MP0/a_216_n18# xb1/MN1/a_324_334#
+ AVSS xb2_1/MN0/a_324_n18# SUNTRB_IVX1_CV
Xxb2_1 AVDD VDD_ROSC AVSS xb2_1/A xb2_2/A xb2_1/MP0/a_216_n18# xb2_2/MP0/a_216_n18#
+ xb2_1/MN0/a_324_n18# AVSS xb2_2/MN0/a_324_n18# SUNTRB_IVX1_CV
C0 xa5/MP0/a_216_n18# AVDD -0.311f
C1 xa6/MP1/a_216_n18# AVDD -0.311f
C2 xb1/B xa3/AN 0.131f
C3 xb2_6/MP0/a_216_n18# AVDD -0.311f
C4 xb2_3/A xb2_4/A 0.134f
C5 xa4/A xa3/AN 0.121f
C6 xb1/B xb1/Y 0.112f
C7 xa4/MP0/a_216_n18# AVDD -0.311f
C8 VDD_ROSC AVDD 0.154f
C9 AVDD xa3/A 0.406f
C10 xb2_5/MP0/a_216_n18# AVDD -0.31f
C11 AVDD xb2_1/MP0/a_216_n18# -0.31f
C12 xb2_3/A xb2_2/A 0.134f
C13 xb2_4/MP0/a_216_n18# AVDD -0.31f
C14 AVDD xa3/AN 0.283f
C15 xb1/MP1/a_216_334# AVDD -0.31f
C16 AVDD xa4/A 0.103f
C17 PWRUP_1V8 AVDD 0.302f
C18 AVDD CK 0.436f
C19 xb2_3/MP0/a_216_n18# AVDD -0.31f
C20 xb2_2/MP0/a_216_n18# AVDD -0.31f
C21 xa5/A xa4/A 0.241f
C22 xb2_5/A xa3/A 0.165f
C23 xb2_2/A xb2_1/A 0.134f
C24 VDD_ROSC xa3/A 0.305f
C25 xb2_1/A xb1/Y 0.121f
C26 xb2_4/A xb2_5/A 0.134f
C27 xa5/A AVDD 0.115f
C28 xb3/MP1/a_216_n18# AVDD -0.311f
C29 VDD_ROSC xa3/AN 0.302f
C30 xa3/AN xa3/A 0.957f
C31 xa4/A xa3/A 0.288f
C32 xb2_7/MP0/a_216_n18# AVDD -0.311f
C33 xb2_1/MN0/a_324_n18# AVSS 0.352f
C34 xb2_1/A AVSS 0.786f
C35 xb1/Y AVSS 0.92f
C36 xa6/MN1/a_324_334# AVSS 0.422f
C37 AVDD AVSS 36.8f
C38 CK AVSS 1.57f
C39 xa5/MN0/a_324_n18# AVSS 0.356f
C40 xa6/MN1/a_324_n18# AVSS 0.354f
C41 xa4/Y AVSS 0.319f
C42 xa4/MN0/a_324_n18# AVSS 0.352f
C43 xa3/xb2_1/a_324_n18# AVSS 0.355f
C44 xa3/A AVSS 3.01f
C45 xa3/xb2_0/a_324_n18# AVSS 0.355f
C46 xa3/xb1_1/a_324_n18# AVSS 0.352f
C47 xa3/AN AVSS 2.99f
C48 xa4/A AVSS 1.57f
C49 xa3/xb1_0/a_324_n18# AVSS 0.467f
C50 xa5/A AVSS 1.15f
C51 xa3/xc1a/a_216_n18# AVSS 0.13f
C52 xb3/MN1/a_324_334# AVSS 0.461f
C53 xb3/MP1/S AVSS 0.233f
C54 xb3/MP1/a_216_334# AVSS 0.129f
C55 xb1/MN1/a_324_334# AVSS 0.353f
C56 VDD_ROSC AVSS 0.785f
C57 xb1/MN0/a_324_n18# AVSS 0.469f
C58 xb1/MN1/a_324_n18# AVSS 0.358f
C59 xb1/B AVSS 2.5f
C60 PWRUP_1V8 AVSS 1.23f
C61 xb1/MP0/a_216_n18# AVSS 0.131f
C62 xb3/MN1/a_324_n18# AVSS 0.354f
C63 xb2_6/MN0/a_324_n18# AVSS 0.349f
C64 xb2_7/MN0/a_324_n18# AVSS 0.349f
C65 xb2_5/MN0/a_324_n18# AVSS 0.352f
C66 xb2_5/A AVSS 0.782f
C67 xb2_4/MN0/a_324_n18# AVSS 0.352f
C68 xb2_4/A AVSS 0.782f
C69 xb2_2/MN0/a_324_n18# AVSS 0.352f
C70 xb2_2/A AVSS 0.782f
C71 xb2_3/MN0/a_324_n18# AVSS 0.352f
C72 xb2_3/A AVSS 0.782f
.ends

.subckt SUNTR_NDX1_CV B Y AVDD AVSS MN1/a_324_334# A MP1/B MP0/a_216_n18# MP1/a_216_334#
+ MN0/a_324_n18# VSUBS
XMP0 Y A AVDD MP1/B MP0/a_216_n18# MP1/a_216_n18# VSUBS SUNTR_PCHDL
XMP1 AVDD B Y MP1/B MP1/a_216_n18# MP1/a_216_334# VSUBS SUNTR_PCHDL
XMN0 MN1/S A AVSS VSUBS MN0/a_324_n18# MN1/a_324_n18# SUNTR_NCHDL
XMN1 Y B MN1/S VSUBS MN1/a_324_n18# MN1/a_324_334# SUNTR_NCHDL
C0 MP1/a_216_n18# MP1/B -0.311f
C1 MP1/B AVDD 0.175f
C2 MP1/B B 0.11f
C3 MP1/B Y 0.115f
C4 MP1/B A 0.11f
C5 AVDD VSUBS 0.345f
C6 AVSS VSUBS 0.411f
C7 B VSUBS 0.561f
C8 Y VSUBS 0.299f
C9 MN1/a_324_n18# VSUBS 0.352f
C10 MN1/a_324_334# VSUBS 0.422f
C11 A VSUBS 0.562f
C12 MN0/a_324_n18# VSUBS 0.422f
C13 MP1/B VSUBS 4.38f
.ends

.subckt SUNTR_IVTRIX1_CV CN AVDD AVSS MN1/a_324_334# C Y MP1/B MP0/a_216_n18# MP1/a_216_334#
+ A MN0/a_324_n18# VSUBS
XMP0 MP1/S A AVDD MP1/B MP0/a_216_n18# MP1/a_216_n18# VSUBS SUNTR_PCHDL
XMP1 Y CN MP1/S MP1/B MP1/a_216_n18# MP1/a_216_334# VSUBS SUNTR_PCHDL
XMN0 MN1/S A AVSS VSUBS MN0/a_324_n18# MN1/a_324_n18# SUNTR_NCHDL
XMN1 Y C MN1/S VSUBS MN1/a_324_n18# MN1/a_324_334# SUNTR_NCHDL
C0 MP1/B AVDD 0.137f
C1 MP1/B A 0.116f
C2 MP1/a_216_n18# MP1/B -0.311f
C3 AVDD VSUBS 0.272f
C4 AVSS VSUBS 0.415f
C5 A VSUBS 0.579f
C6 C VSUBS 0.384f
C7 Y VSUBS 0.255f
C8 MN1/a_324_n18# VSUBS 0.352f
C9 MN1/a_324_334# VSUBS 0.422f
C10 MN0/a_324_n18# VSUBS 0.422f
C11 MP1/B VSUBS 4.38f
.ends

.subckt SUNTR_NDTRIX1_CV C CN Y AVDD AVSS MN1/a_324_334# MN2/a_324_n18# MP2/B RN MP2/S
+ MP1/a_216_334# A MP2/a_216_n18# VSUBS
XMP0 MP2/S A AVDD MP2/B MP2/a_216_334# MP1/a_216_n18# VSUBS SUNTR_PCHDL
XMP1 Y CN MP2/S MP2/B MP1/a_216_n18# MP1/a_216_334# VSUBS SUNTR_PCHDL
XMP2 AVDD RN MP2/S MP2/B MP2/a_216_n18# MP2/a_216_334# VSUBS SUNTR_PCHDL
XMN0 MP2/S A MN2/D VSUBS MN2/a_324_334# MN1/a_324_n18# SUNTR_NCHDL
XMN1 Y C MP2/S VSUBS MN1/a_324_n18# MN1/a_324_334# SUNTR_NCHDL
XMN2 MN2/D RN AVSS VSUBS MN2/a_324_n18# MN2/a_324_334# SUNTR_NCHDL
C0 MP2/B AVDD 0.18f
C1 MP2/B A 0.116f
C2 MP2/B RN 0.109f
C3 MP2/B MP2/S 0.188f
C4 MP2/B MP2/a_216_334# -0.311f
C5 AVSS AVDD 0.12f
C6 MP1/a_216_n18# MP2/B -0.311f
C7 MP2/S AVDD 0.161f
C8 AVDD VSUBS 0.301f
C9 A VSUBS 0.512f
C10 AVSS VSUBS 0.484f
C11 RN VSUBS 0.562f
C12 MN2/a_324_n18# VSUBS 0.422f
C13 MN2/a_324_334# VSUBS 0.352f
C14 C VSUBS 0.384f
C15 Y VSUBS 0.216f
C16 MN1/a_324_n18# VSUBS 0.352f
C17 MN1/a_324_334# VSUBS 0.422f
C18 MP2/S VSUBS 0.252f
C19 MP2/B VSUBS 5.96f
.ends

.subckt SUNTR_DFRNQNX1_CV RN Q XA5/A D QN XA7/C XA6/A CK AVDD AVSS
XXA0 AVDD XA0/MN1/a_324_n18# XA1/MN0/a_324_n18# XA1/MP0/a_216_n18# XA0/MP1/a_216_n18#
+ AVSS SUNTR_TAPCELLB_CV
XXA1 RN XA7/C AVDD AVSS XA2/MN0/a_324_n18# CK AVDD XA1/MP0/a_216_n18# XA2/MP0/a_216_n18#
+ XA1/MN0/a_324_n18# AVSS SUNTR_NDX1_CV
XXA2 AVDD AVSS AVDD XA6/C XA2/MP0/a_216_n18# XA3/MP0/a_216_n18# XA7/C XA2/MN0/a_324_n18#
+ AVSS XA3/MN0/a_324_n18# SUNTR_IVX1_CV
XXA3 XA6/C AVDD AVSS XA4/MN0/a_324_n18# XA7/C XA5/A AVDD XA3/MP0/a_216_n18# XA4/MP0/a_216_n18#
+ D XA3/MN0/a_324_n18# AVSS SUNTR_IVTRIX1_CV
XXA5 AVDD AVSS AVDD XA6/A XA5/MP0/a_216_n18# XA6/MP0/a_216_n18# XA5/A XA5/MN0/a_324_n18#
+ AVSS XA6/MN0/a_324_n18# SUNTR_IVX1_CV
XXA4 XA7/C AVDD AVSS XA5/MN0/a_324_n18# XA6/C XA5/A AVDD XA4/MP0/a_216_n18# XA5/MP0/a_216_n18#
+ XA6/A XA4/MN0/a_324_n18# AVSS SUNTR_IVTRIX1_CV
XXA6 XA7/C AVDD AVSS XA7/MN2/a_324_n18# XA6/C QN AVDD XA6/MP0/a_216_n18# XA7/MP2/a_216_n18#
+ XA6/A XA6/MN0/a_324_n18# AVSS SUNTR_IVTRIX1_CV
XXA7 XA7/C XA6/C QN AVDD AVSS XA8/MN0/a_324_n18# XA7/MN2/a_324_n18# AVDD RN XA7/MP2/S
+ XA8/MP0/a_216_n18# Q XA7/MP2/a_216_n18# AVSS SUNTR_NDTRIX1_CV
XXA8 AVDD AVSS AVDD Q XA8/MP0/a_216_n18# XA8/MP0/a_216_334# QN XA8/MN0/a_324_n18#
+ AVSS XA8/MN0/a_324_334# SUNTR_IVX1_CV
C0 XA7/C QN 0.157f
C1 XA6/C XA7/MP2/S 0.107f
C2 AVSS QN 0.392f
C3 AVDD XA8/MP0/a_216_n18# -0.312f
C4 XA7/C RN 0.379f
C5 XA6/C RN 0.116f
C6 AVDD QN 0.151f
C7 AVSS RN 0.436f
C8 QN Q 0.162f
C9 AVDD XA3/MP0/a_216_n18# -0.313f
C10 XA7/C XA6/A 0.294f
C11 XA6/C XA6/A 0.489f
C12 AVDD XA7/MP2/a_216_n18# -0.314f
C13 XA6/C XA7/C 0.465f
C14 AVSS XA7/C 0.678f
C15 AVSS XA6/C 0.275f
C16 XA5/A XA6/A 0.216f
C17 XA6/C XA5/A 0.367f
C18 AVSS XA5/A 0.272f
C19 AVDD XA6/A 0.558f
C20 AVDD XA7/C 1.99f
C21 AVDD XA6/C 1.17f
C22 QN XA7/MP2/S 0.193f
C23 XA6/C Q 0.174f
C24 AVDD XA5/A 0.164f
C25 AVDD XA6/MP0/a_216_n18# -0.315f
C26 AVDD XA2/MP0/a_216_n18# -0.313f
C27 XA6/C D 0.101f
C28 XA1/MP0/a_216_n18# AVDD -0.312f
C29 AVDD Q 0.371f
C30 XA5/MP0/a_216_n18# AVDD -0.313f
C31 AVDD XA4/MP0/a_216_n18# -0.313f
C32 QN 0 1.18f
C33 Q 0 0.85f
C34 XA8/MN0/a_324_n18# 0 0.36f
C35 XA8/MN0/a_324_334# 0 0.422f
C36 XA7/MN2/a_324_n18# 0 0.36f
C37 XA7/MN2/a_324_334# 0 0.355f
C38 XA7/MN1/a_324_n18# 0 0.355f
C39 XA7/MP2/S 0 0.246f
C40 XA6/MN1/a_324_n18# 0 0.355f
C41 XA6/MN0/a_324_n18# 0 0.36f
C42 XA6/A 0 1.13f
C43 XA5/A 0 0.931f
C44 XA4/MN1/a_324_n18# 0 0.355f
C45 XA4/MN0/a_324_n18# 0 0.36f
C46 XA5/MN0/a_324_n18# 0 0.36f
C47 D 0 0.499f
C48 XA3/MN1/a_324_n18# 0 0.355f
C49 XA3/MN0/a_324_n18# 0 0.36f
C50 XA7/C 0 2.72f
C51 XA6/C 0 1.47f
C52 RN 0 2.04f
C53 XA1/MN1/a_324_n18# 0 0.355f
C54 XA2/MN0/a_324_n18# 0 0.36f
C55 CK 0 0.512f
C56 XA1/MN0/a_324_n18# 0 0.36f
C57 AVSS 0 0.147f
C58 XA0/MN1/a_324_n18# 0 0.422f
C59 AVDD 0 25.3f
.ends

.subckt SUN_PLL_DIVN CK_FB CK PWRUP_1V8 AVDD AVSS
Xxc PWRUP_1V8 CK_FB xc/XA5/A xc/D xc/D xc/XA7/C xc/XA6/A xd/Q AVDD AVSS SUNTR_DFRNQNX1_CV
Xxd PWRUP_1V8 xd/Q xd/XA5/A xd/D xd/D xd/XA7/C xd/XA6/A xe/Q AVDD AVSS SUNTR_DFRNQNX1_CV
Xxe PWRUP_1V8 xe/Q xe/XA5/A xe/D xe/D xe/XA7/C xe/XA6/A xf/Q AVDD AVSS SUNTR_DFRNQNX1_CV
Xxf PWRUP_1V8 xf/Q xf/XA5/A xf/D xf/D xf/XA7/C xf/XA6/A xg/Q AVDD AVSS SUNTR_DFRNQNX1_CV
Xxg PWRUP_1V8 xg/Q xg/XA5/A xg/D xg/D xg/XA7/C xg/XA6/A CK AVDD AVSS SUNTR_DFRNQNX1_CV
C0 xf/Q AVSS 0.729f
C1 xe/XA6/C xe/D 0.109f
C2 AVDD CK_FB 0.245f
C3 xd/XA7/C xd/Q 0.146f
C4 xg/XA6/A xg/D 0.185f
C5 xf/XA7/C xf/Q 0.146f
C6 PWRUP_1V8 xg/Q 0.41f
C7 xe/Q PWRUP_1V8 0.41f
C8 xf/Q AVDD 1.99f
C9 xd/XA7/C xc/XA7/C 0.31f
C10 xc/D xc/XA6/A 0.185f
C11 xf/XA7/C xe/XA7/C 0.31f
C12 xc/XA7/C xc/D 0.161f
C13 xc/XA6/C xc/D 0.109f
C14 xe/XA6/A xe/D 0.185f
C15 AVSS xc/D 0.264f
C16 xc/D xc/XA5/A 0.286f
C17 xg/XA7/C xg/Q 0.14f
C18 xg/XA7/C PWRUP_1V8 0.182f
C19 xc/XA7/C PWRUP_1V8 0.191f
C20 xe/XA5/A xe/D 0.286f
C21 AVDD xc/D 0.512f
C22 xd/D xd/XA6/A 0.185f
C23 AVSS xg/Q 1.08f
C24 xe/Q AVSS 1.07f
C25 AVSS PWRUP_1V8 2.07f
C26 xd/XA7/C xd/D 0.161f
C27 xe/XA7/C xf/Q 0.298f
C28 xd/XA6/C xd/D 0.109f
C29 xd/Q xc/XA7/C 0.298f
C30 xf/XA7/C xg/Q 0.11f
C31 xf/XA7/C PWRUP_1V8 0.191f
C32 xd/Q AVSS 0.734f
C33 xg/XA5/A xg/D 0.286f
C34 xd/D xd/XA5/A 0.286f
C35 xe/Q AVDD 0.111f
C36 AVDD PWRUP_1V8 2.62f
C37 AVSS xg/XA7/C 0.101f
C38 xg/XA7/C xg/D 0.161f
C39 xe/D AVSS 0.262f
C40 AVSS CK 0.401f
C41 PWRUP_1V8 CK_FB 0.162f
C42 xd/Q AVDD 1.99f
C43 AVSS xg/D 0.263f
C44 xg/XA6/C xg/D 0.109f
C45 xe/D AVDD 0.512f
C46 xf/XA6/A xf/D 0.185f
C47 AVDD CK 0.308f
C48 xe/XA7/C xe/Q 0.14f
C49 xe/XA7/C PWRUP_1V8 0.182f
C50 AVDD AVSS 11.2f
C51 AVDD xg/D 0.508f
C52 xd/D AVSS 0.262f
C53 xf/D AVSS 0.262f
C54 AVSS CK_FB 0.408f
C55 xf/XA5/A xf/D 0.286f
C56 xf/XA7/C xf/D 0.161f
C57 xd/XA7/C xe/Q 0.11f
C58 xd/XA7/C PWRUP_1V8 0.191f
C59 xf/XA6/C xf/D 0.109f
C60 xd/D AVDD 0.512f
C61 xf/D AVDD 0.512f
C62 xe/XA7/C xe/D 0.161f
C63 xg/D 0 1.93f
C64 xg/Q 0 2.37f
C65 xg/XA8/MN0/a_324_n18# 0 0.36f
C66 xg/XA8/MN0/a_324_334# 0 0.422f
C67 xg/XA7/MN2/a_324_n18# 0 0.36f
C68 xg/XA7/MN2/a_324_334# 0 0.355f
C69 xg/XA7/MN1/a_324_n18# 0 0.355f
C70 xg/XA7/MP2/S 0 0.246f
C71 xg/XA6/MN1/a_324_n18# 0 0.355f
C72 xg/XA6/MN0/a_324_n18# 0 0.36f
C73 xg/XA6/A 0 1.13f
C74 xg/XA5/A 0 0.931f
C75 xg/XA4/MN1/a_324_n18# 0 0.355f
C76 xg/XA4/MN0/a_324_n18# 0 0.36f
C77 xg/XA5/MN0/a_324_n18# 0 0.36f
C78 xg/XA3/MN1/a_324_n18# 0 0.355f
C79 xg/XA3/MN0/a_324_n18# 0 0.36f
C80 xg/XA7/C 0 2.72f
C81 xg/XA6/C 0 1.47f
C82 xg/XA1/MN1/a_324_n18# 0 0.355f
C83 xg/XA2/MN0/a_324_n18# 0 0.36f
C84 CK 0 0.934f
C85 xg/XA1/MN0/a_324_n18# 0 0.36f
C86 xg/XA0/MN1/a_324_n18# 0 0.422f
C87 xf/D 0 1.92f
C88 xf/Q 0 2.11f
C89 xf/XA8/MN0/a_324_n18# 0 0.36f
C90 xf/XA8/MN0/a_324_334# 0 0.422f
C91 xf/XA7/MN2/a_324_n18# 0 0.36f
C92 xf/XA7/MN2/a_324_334# 0 0.355f
C93 xf/XA7/MN1/a_324_n18# 0 0.355f
C94 xf/XA7/MP2/S 0 0.246f
C95 xf/XA6/MN1/a_324_n18# 0 0.355f
C96 xf/XA6/MN0/a_324_n18# 0 0.36f
C97 xf/XA6/A 0 1.13f
C98 xf/XA5/A 0 0.931f
C99 xf/XA4/MN1/a_324_n18# 0 0.355f
C100 xf/XA4/MN0/a_324_n18# 0 0.36f
C101 xf/XA5/MN0/a_324_n18# 0 0.36f
C102 xf/XA3/MN1/a_324_n18# 0 0.355f
C103 xf/XA3/MN0/a_324_n18# 0 0.36f
C104 xf/XA7/C 0 2.72f
C105 xf/XA6/C 0 1.47f
C106 xf/XA1/MN1/a_324_n18# 0 0.355f
C107 xf/XA2/MN0/a_324_n18# 0 0.36f
C108 xf/XA1/MN0/a_324_n18# 0 0.36f
C109 xf/XA0/MN1/a_324_n18# 0 0.422f
C110 xe/D 0 1.93f
C111 xe/Q 0 2.32f
C112 xe/XA8/MN0/a_324_n18# 0 0.36f
C113 xe/XA8/MN0/a_324_334# 0 0.422f
C114 xe/XA7/MN2/a_324_n18# 0 0.36f
C115 xe/XA7/MN2/a_324_334# 0 0.355f
C116 xe/XA7/MN1/a_324_n18# 0 0.355f
C117 xe/XA7/MP2/S 0 0.246f
C118 xe/XA6/MN1/a_324_n18# 0 0.355f
C119 xe/XA6/MN0/a_324_n18# 0 0.36f
C120 xe/XA6/A 0 1.13f
C121 xe/XA5/A 0 0.931f
C122 xe/XA4/MN1/a_324_n18# 0 0.355f
C123 xe/XA4/MN0/a_324_n18# 0 0.36f
C124 xe/XA5/MN0/a_324_n18# 0 0.36f
C125 xe/XA3/MN1/a_324_n18# 0 0.355f
C126 xe/XA3/MN0/a_324_n18# 0 0.36f
C127 xe/XA7/C 0 2.72f
C128 xe/XA6/C 0 1.47f
C129 xe/XA1/MN1/a_324_n18# 0 0.355f
C130 xe/XA2/MN0/a_324_n18# 0 0.36f
C131 xe/XA1/MN0/a_324_n18# 0 0.36f
C132 xe/XA0/MN1/a_324_n18# 0 0.422f
C133 xd/D 0 1.92f
C134 xd/Q 0 2.13f
C135 xd/XA8/MN0/a_324_n18# 0 0.36f
C136 xd/XA8/MN0/a_324_334# 0 0.422f
C137 xd/XA7/MN2/a_324_n18# 0 0.36f
C138 xd/XA7/MN2/a_324_334# 0 0.355f
C139 xd/XA7/MN1/a_324_n18# 0 0.355f
C140 xd/XA7/MP2/S 0 0.246f
C141 xd/XA6/MN1/a_324_n18# 0 0.355f
C142 xd/XA6/MN0/a_324_n18# 0 0.36f
C143 xd/XA6/A 0 1.13f
C144 xd/XA5/A 0 0.931f
C145 xd/XA4/MN1/a_324_n18# 0 0.355f
C146 xd/XA4/MN0/a_324_n18# 0 0.36f
C147 xd/XA5/MN0/a_324_n18# 0 0.36f
C148 xd/XA3/MN1/a_324_n18# 0 0.355f
C149 xd/XA3/MN0/a_324_n18# 0 0.36f
C150 xd/XA7/C 0 2.72f
C151 xd/XA6/C 0 1.47f
C152 xd/XA1/MN1/a_324_n18# 0 0.355f
C153 xd/XA2/MN0/a_324_n18# 0 0.36f
C154 xd/XA1/MN0/a_324_n18# 0 0.36f
C155 xd/XA0/MN1/a_324_n18# 0 0.422f
C156 xc/D 0 1.93f
C157 CK_FB 0 1.02f
C158 xc/XA8/MN0/a_324_n18# 0 0.36f
C159 xc/XA8/MN0/a_324_334# 0 0.422f
C160 xc/XA7/MN2/a_324_n18# 0 0.36f
C161 xc/XA7/MN2/a_324_334# 0 0.355f
C162 xc/XA7/MN1/a_324_n18# 0 0.355f
C163 xc/XA7/MP2/S 0 0.246f
C164 xc/XA6/MN1/a_324_n18# 0 0.355f
C165 xc/XA6/MN0/a_324_n18# 0 0.36f
C166 xc/XA6/A 0 1.13f
C167 xc/XA5/A 0 0.931f
C168 xc/XA4/MN1/a_324_n18# 0 0.355f
C169 xc/XA4/MN0/a_324_n18# 0 0.36f
C170 xc/XA5/MN0/a_324_n18# 0 0.36f
C171 xc/XA3/MN1/a_324_n18# 0 0.355f
C172 xc/XA3/MN0/a_324_n18# 0 0.36f
C173 xc/XA7/C 0 2.72f
C174 xc/XA6/C 0 1.47f
C175 PWRUP_1V8 0 17f
C176 xc/XA1/MN1/a_324_n18# 0 0.355f
C177 xc/XA2/MN0/a_324_n18# 0 0.36f
C178 xc/XA1/MN0/a_324_n18# 0 0.36f
C179 AVSS 0 -3.74f
C180 xc/XA0/MN1/a_324_n18# 0 0.422f
C181 AVDD 0 0.117p
.ends

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt SUN_PLL AVDD AVSS PWRUP_1V8 CK_REF CK IBPSR_1U
*.subckt SUN_PLL AVDD AVSS PWRUP_1V8 CK_REF CK IBPSR_1U
Xxbb1 IBPSR_1U xbb1/PWRUP_1V8_N AVSS SUN_PLL_BIAS
Xxbb0 VLPZ VLPF AVSS SUN_PLL_LPF
Xxaa0 xaa1/CP_UP_N CK_REF xaa1/CP_DOWN xaa6/CK_FB AVDD xaa0/xa5/D AVSS SUN_PLL_PFD
Xxaa1 AVDD xaa1/CP_UP_N VLPF xaa1/CP_DOWN IBPSR_1U VLPZ PWRUP_1V8 xaa3/KICK AVSS SUN_PLL_CP
Xxaa3 xaa3/KICK xaa3/KICK_N xbb1/PWRUP_1V8_N AVDD AVSS PWRUP_1V8 SUN_PLL_KICK
Xxaa4 AVDD VDD_ROSC VLPF VDD_ROSC IBPSR_1U AVSS SUN_PLL_BUF
Xxaa5 AVDD CK VDD_ROSC PWRUP_1V8 AVSS SUN_PLL_ROSC
Xxaa6 xaa6/CK_FB CK PWRUP_1V8 AVDD AVSS SUN_PLL_DIVN
C0 xbb0/xa2/N VLPZ 0.448f
C1 AVDD xaa6/CK_FB 2.35f
C2 xaa1/CP_DOWN AVDD 0.641f
C3 VDD_ROSC AVSS 0.749f
C4 VLPZ AVSS 0.871f
C5 xaa3/KICK AVDD 1.61f
C6 CK PWRUP_1V8 0.21f
C7 xbb1/PWRUP_1V8_N IBPSR_1U 0.765f
C8 VDD_ROSC AVDD 2.66f
C9 VLPF VDD_ROSC 0.1f
C10 VLPZ AVDD 0.776f
C11 VLPF VLPZ 3.39f
C12 xbb0/xa1/XA1/a_n72_n110# VLPZ 0.181f
C13 IBPSR_1U AVSS 1.85f
C14 xbb1/PWRUP_1V8_N PWRUP_1V8 1.56f
C15 xaa1/CP_UP_N AVDD 0.265f
C16 AVSS PWRUP_1V8 6.98f
C17 xaa3/KICK VLPZ 0.181f
C18 IBPSR_1U AVDD 1.56f
C19 CK AVSS 2.9f
C20 PWRUP_1V8 xaa0/xa5/D 0.238f
C21 xaa1/CP_UP_N xaa1/CP_DOWN 3.25f
C22 xaa1/CP_DOWN IBPSR_1U 0.189f
C23 AVDD PWRUP_1V8 6.06f
C24 CK AVDD 2.53f
C25 xbb1/PWRUP_1V8_N AVSS 0.323f
C26 xaa6/xg/XA7/C CK 0.248f
C27 PWRUP_1V8 xaa6/CK_FB 5.18f
C28 xaa1/CP_DOWN PWRUP_1V8 0.181f
C29 xbb1/PWRUP_1V8_N AVDD 0.152f
C30 xaa1/CP_UP_N IBPSR_1U 0.441f
C31 AVDD AVSS 6.63f
C32 VDD_ROSC CK 0.794f
C33 VLPF AVSS 1.53f
C34 AVSS xaa6/CK_FB 5.52f
C35 xbb0/xa2/XA1/a_n72_n110# VLPZ 0.187f
C36 xaa1/CP_DOWN AVSS 0.3f
C37 xaa1/CP_UP_N PWRUP_1V8 0.1f
C38 VLPF AVDD 8.01f
C39 xaa3/KICK AVSS 0.307f
C40 IBPSR_1U PWRUP_1V8 2.33f
C41 xaa6/xg/D 0 1.93f
C42 xaa6/xg/Q 0 2.37f
C43 xaa6/xg/XA8/MN0/a_324_n18# 0 0.36f
C44 xaa6/xg/XA8/MN0/a_324_334# 0 0.422f
C45 xaa6/xg/XA7/MN2/a_324_n18# 0 0.36f
C46 xaa6/xg/XA7/MN2/a_324_334# 0 0.355f
C47 xaa6/xg/XA7/MN1/a_324_n18# 0 0.355f
C48 xaa6/xg/XA7/MP2/S 0 0.246f
C49 xaa6/xg/XA6/MN1/a_324_n18# 0 0.355f
C50 xaa6/xg/XA6/MN0/a_324_n18# 0 0.36f
C51 xaa6/xg/XA6/A 0 1.13f
C52 xaa6/xg/XA5/A 0 0.931f
C53 xaa6/xg/XA4/MN1/a_324_n18# 0 0.355f
C54 xaa6/xg/XA4/MN0/a_324_n18# 0 0.36f
C55 xaa6/xg/XA5/MN0/a_324_n18# 0 0.36f
C56 xaa6/xg/XA3/MN1/a_324_n18# 0 0.355f
C57 xaa6/xg/XA3/MN0/a_324_n18# 0 0.36f
C58 xaa6/xg/XA7/C 0 2.72f
C59 xaa6/xg/XA6/C 0 1.47f
C60 xaa6/xg/XA1/MN1/a_324_n18# 0 0.355f
C61 xaa6/xg/XA2/MN0/a_324_n18# 0 0.36f
C62 CK 0 2.8f
C63 xaa6/xg/XA1/MN0/a_324_n18# 0 0.36f
C64 xaa6/xg/XA0/MN1/a_324_n18# 0 0.422f
C65 xaa6/xf/D 0 1.92f
C66 xaa6/xf/Q 0 2.11f
C67 xaa6/xf/XA8/MN0/a_324_n18# 0 0.36f
C68 xaa6/xf/XA8/MN0/a_324_334# 0 0.422f
C69 xaa6/xf/XA7/MN2/a_324_n18# 0 0.36f
C70 xaa6/xf/XA7/MN2/a_324_334# 0 0.355f
C71 xaa6/xf/XA7/MN1/a_324_n18# 0 0.355f
C72 xaa6/xf/XA7/MP2/S 0 0.246f
C73 xaa6/xf/XA6/MN1/a_324_n18# 0 0.355f
C74 xaa6/xf/XA6/MN0/a_324_n18# 0 0.36f
C75 xaa6/xf/XA6/A 0 1.13f
C76 xaa6/xf/XA5/A 0 0.931f
C77 xaa6/xf/XA4/MN1/a_324_n18# 0 0.355f
C78 xaa6/xf/XA4/MN0/a_324_n18# 0 0.36f
C79 xaa6/xf/XA5/MN0/a_324_n18# 0 0.36f
C80 xaa6/xf/XA3/MN1/a_324_n18# 0 0.355f
C81 xaa6/xf/XA3/MN0/a_324_n18# 0 0.36f
C82 xaa6/xf/XA7/C 0 2.72f
C83 xaa6/xf/XA6/C 0 1.47f
C84 xaa6/xf/XA1/MN1/a_324_n18# 0 0.355f
C85 xaa6/xf/XA2/MN0/a_324_n18# 0 0.36f
C86 xaa6/xf/XA1/MN0/a_324_n18# 0 0.36f
C87 xaa6/xf/XA0/MN1/a_324_n18# 0 0.422f
C88 xaa6/xe/D 0 1.93f
C89 xaa6/xe/Q 0 2.32f
C90 xaa6/xe/XA8/MN0/a_324_n18# 0 0.36f
C91 xaa6/xe/XA8/MN0/a_324_334# 0 0.422f
C92 xaa6/xe/XA7/MN2/a_324_n18# 0 0.36f
C93 xaa6/xe/XA7/MN2/a_324_334# 0 0.355f
C94 xaa6/xe/XA7/MN1/a_324_n18# 0 0.355f
C95 xaa6/xe/XA7/MP2/S 0 0.246f
C96 xaa6/xe/XA6/MN1/a_324_n18# 0 0.355f
C97 xaa6/xe/XA6/MN0/a_324_n18# 0 0.36f
C98 xaa6/xe/XA6/A 0 1.13f
C99 xaa6/xe/XA5/A 0 0.931f
C100 xaa6/xe/XA4/MN1/a_324_n18# 0 0.355f
C101 xaa6/xe/XA4/MN0/a_324_n18# 0 0.36f
C102 xaa6/xe/XA5/MN0/a_324_n18# 0 0.36f
C103 xaa6/xe/XA3/MN1/a_324_n18# 0 0.355f
C104 xaa6/xe/XA3/MN0/a_324_n18# 0 0.36f
C105 xaa6/xe/XA7/C 0 2.72f
C106 xaa6/xe/XA6/C 0 1.47f
C107 xaa6/xe/XA1/MN1/a_324_n18# 0 0.355f
C108 xaa6/xe/XA2/MN0/a_324_n18# 0 0.36f
C109 xaa6/xe/XA1/MN0/a_324_n18# 0 0.36f
C110 xaa6/xe/XA0/MN1/a_324_n18# 0 0.422f
C111 xaa6/xd/D 0 1.92f
C112 xaa6/xd/Q 0 2.13f
C113 xaa6/xd/XA8/MN0/a_324_n18# 0 0.36f
C114 xaa6/xd/XA8/MN0/a_324_334# 0 0.422f
C115 xaa6/xd/XA7/MN2/a_324_n18# 0 0.36f
C116 xaa6/xd/XA7/MN2/a_324_334# 0 0.355f
C117 xaa6/xd/XA7/MN1/a_324_n18# 0 0.355f
C118 xaa6/xd/XA7/MP2/S 0 0.246f
C119 xaa6/xd/XA6/MN1/a_324_n18# 0 0.355f
C120 xaa6/xd/XA6/MN0/a_324_n18# 0 0.36f
C121 xaa6/xd/XA6/A 0 1.13f
C122 xaa6/xd/XA5/A 0 0.931f
C123 xaa6/xd/XA4/MN1/a_324_n18# 0 0.355f
C124 xaa6/xd/XA4/MN0/a_324_n18# 0 0.36f
C125 xaa6/xd/XA5/MN0/a_324_n18# 0 0.36f
C126 xaa6/xd/XA3/MN1/a_324_n18# 0 0.355f
C127 xaa6/xd/XA3/MN0/a_324_n18# 0 0.36f
C128 xaa6/xd/XA7/C 0 2.72f
C129 xaa6/xd/XA6/C 0 1.47f
C130 xaa6/xd/XA1/MN1/a_324_n18# 0 0.355f
C131 xaa6/xd/XA2/MN0/a_324_n18# 0 0.36f
C132 xaa6/xd/XA1/MN0/a_324_n18# 0 0.36f
C133 xaa6/xd/XA0/MN1/a_324_n18# 0 0.422f
C134 xaa6/xc/D 0 1.93f
C135 xaa6/CK_FB 0 8.86f
C136 xaa6/xc/XA8/MN0/a_324_n18# 0 0.36f
C137 xaa6/xc/XA8/MN0/a_324_334# 0 0.422f
C138 xaa6/xc/XA7/MN2/a_324_n18# 0 0.36f
C139 xaa6/xc/XA7/MN2/a_324_334# 0 0.355f
C140 xaa6/xc/XA7/MN1/a_324_n18# 0 0.355f
C141 xaa6/xc/XA7/MP2/S 0 0.246f
C142 xaa6/xc/XA6/MN1/a_324_n18# 0 0.355f
C143 xaa6/xc/XA6/MN0/a_324_n18# 0 0.36f
C144 xaa6/xc/XA6/A 0 1.13f
C145 xaa6/xc/XA5/A 0 0.931f
C146 xaa6/xc/XA4/MN1/a_324_n18# 0 0.355f
C147 xaa6/xc/XA4/MN0/a_324_n18# 0 0.36f
C148 xaa6/xc/XA5/MN0/a_324_n18# 0 0.36f
C149 xaa6/xc/XA3/MN1/a_324_n18# 0 0.355f
C150 xaa6/xc/XA3/MN0/a_324_n18# 0 0.36f
C151 xaa6/xc/XA7/C 0 2.72f
C152 xaa6/xc/XA6/C 0 1.47f
C153 PWRUP_1V8 0 27.9f
C154 xaa6/xc/XA1/MN1/a_324_n18# 0 0.355f
C155 xaa6/xc/XA2/MN0/a_324_n18# 0 0.36f
C156 xaa6/xc/XA1/MN0/a_324_n18# 0 0.36f
C157 AVSS 0 1.38p
C158 xaa6/xc/XA0/MN1/a_324_n18# 0 0.422f
C159 AVDD 0 0.298p
C160 xaa5/xb2_1/MN0/a_324_n18# 0 0.36f
C161 xaa5/xb2_1/A 0 0.669f
C162 xaa5/xb1/Y 0 0.764f
C163 xaa5/xa6/MN1/a_324_334# 0 0.422f
C164 xaa5/xa5/MN0/a_324_n18# 0 0.36f
C165 xaa5/xa6/MN1/a_324_n18# 0 0.36f
C166 xaa5/xa4/Y 0 0.264f
C167 xaa5/xa4/MN0/a_324_n18# 0 0.36f
C168 xaa5/xa3/xb2_1/a_324_n18# 0 0.355f
C169 xaa5/xa3/A 0 2.15f
C170 xaa5/xa3/xb2_0/a_324_n18# 0 0.355f
C171 xaa5/xa3/xb1_1/a_324_n18# 0 0.355f
C172 xaa5/xa3/AN 0 2.15f
C173 xaa5/xa4/A 0 1.2f
C174 xaa5/xa3/xb1_0/a_324_n18# 0 0.422f
C175 xaa5/xa5/A 0 0.922f
C176 xaa5/xb3/MN1/a_324_334# 0 0.422f
C177 xaa5/xb3/MP1/S 0 0.177f
C178 xaa5/xb1/MN1/a_324_334# 0 0.36f
C179 xaa5/xb1/MN0/a_324_n18# 0 0.422f
C180 xaa5/xb1/MN1/a_324_n18# 0 0.355f
C181 xaa5/xb1/B 0 1.29f
C182 xaa5/xb3/MN1/a_324_n18# 0 0.36f
C183 xaa5/xb2_6/MN0/a_324_n18# 0 0.36f
C184 xaa5/xb2_7/MN0/a_324_n18# 0 0.36f
C185 xaa5/xb2_5/MN0/a_324_n18# 0 0.36f
C186 xaa5/xb2_5/A 0 0.668f
C187 xaa5/xb2_4/MN0/a_324_n18# 0 0.36f
C188 xaa5/xb2_4/A 0 0.665f
C189 xaa5/xb2_2/MN0/a_324_n18# 0 0.36f
C190 xaa5/xb2_2/A 0 0.665f
C191 xaa5/xb2_3/MN0/a_324_n18# 0 0.36f
C192 xaa5/xb2_3/A 0 0.665f
C193 xaa4/xc2_3/G 0 1.59f
C194 xaa4/xc3_9/G 0 2.04f
C195 xaa4/xc3_9/a_216_492# 0 0.106f
C196 xaa4/xc1_0/a_216_n36# 0 0.106f
C197 xaa4/xa4_0/M0/a_324_n18# 0 0.357f
C198 xaa4/xa2_1/M0/a_324_n18# 0 0.357f
C199 VDD_ROSC 0 0.153p
C200 xaa4/xa1/M8/a_324_334# 0 0.357f
C201 xaa4/xa4_1/M8/a_324_334# 0 0.422f
C202 xaa4/xa4_1/M0/a_324_n18# 0 0.357f
C203 VLPF 0 0.157p
C204 xaa4/xa1/D 0 1.44f
C205 xaa4/xa1/M0/a_324_n18# 0 0.422f
C206 xaa3/xa9/MN0/a_324_334# 0 0.422f
C207 xaa3/KICK 0 4.01f
C208 xaa3/xa8/MN1/a_324_n18# 0 0.355f
C209 xaa3/xa9/MN0/a_324_n18# 0 0.36f
C210 xaa3/xa8/MN0/a_324_n18# 0 0.36f
C211 xaa3/xa8/B 0 0.768f
C212 xaa3/xa7/MN0/a_324_n18# 0 0.36f
C213 xaa3/xa7/A 0 0.716f
C214 xaa3/xa6/MN0/a_324_n18# 0 0.422f
C215 xaa3/xa2/MN0/a_324_n18# 0 0.36f
C216 xaa3/xa2/A 0 0.703f
C217 xaa3/xa1c/MN0/a_324_n18# 0 0.36f
C218 xbb1/PWRUP_1V8_N 0 3.5f
C219 xaa3/xa1b/MN0/a_324_n18# 0 0.36f
C220 xaa3/xa1a/MN1/a_324_n18# 0 0.422f
C221 xaa3/xa2/Y 0 0.756f
C222 xaa3/xa6/A 0 2.53f
C223 xaa3/xa2/MN0/a_324_334# 0 0.36f
C224 xaa3/xa5a/MN0/a_324_334# 0 0.422f
C225 xaa1/xa4/M1/a_324_334# 0 0.422f
C226 xaa1/xa3/a_324_334# 0 0.358f
C227 xaa1/xa3/S 0 0.114f
C228 xaa1/xa3/a_324_n18# 0 0.358f
C229 xaa1/xa2/M0/a_324_n18# 0 0.356f
C230 xaa1/xa1/M0/a_324_n18# 0 0.422f
C231 xaa1/xb2/G 0 0.552f
C232 xaa1/CP_DOWN 0 2.61f
C233 xaa0/xa6/MN0/a_324_n18# 0 0.36f
C234 xaa0/xa6/MN0/a_324_334# 0 0.422f
C235 xaa0/xa5/MN2/a_324_n18# 0 0.355f
C236 xaa0/xa5/MN2/a_324_334# 0 0.355f
C237 xaa0/xa5/MP2/G 0 1.03f
C238 xaa0/xa5/MN0/a_324_n18# 0 0.36f
C239 xaa0/xa6/A 0 1.62f
C240 xaa0/xa3/MN1/a_324_n18# 0 0.355f
C241 xaa0/xa3/MN0/a_324_n18# 0 0.36f
C242 xaa0/xa3/A 0 1.5f
C243 xaa0/xa2/MN0/a_324_n18# 0 0.36f
C244 xaa0/xa2/MN0/a_324_334# 0 0.36f
C245 CK_REF 0 0.8f
C246 xaa0/xa1/MN2/a_324_n18# 0 0.355f
C247 xaa0/xa1/MN2/a_324_334# 0 0.355f
C248 xaa0/xa5/D 0 1.97f
C249 xaa0/xa1/MP2/G 0 1.03f
C250 xaa0/xa1/MN0/a_324_n18# 0 0.36f
C251 xaa0/xa0/MN1/a_324_n18# 0 0.422f
C252 xaa0/xa2/Y 0 0.716f
C253 xaa1/CP_UP_N 0 2.43f
C254 VLPZ 0 1.04p
C255 xbb0/xa2/XA1/a_3816_n110# 0 2.55f
C256 xbb0/xa2/XA1/a_2952_n110# 0 0.893f $ **FLOATING
C257 xbb0/xa2/XA1/a_2520_2090# 0 1.1f $ **FLOATING
C258 xbb0/xa2/XA1/a_2088_n110# 0 0.807f $ **FLOATING
C259 xbb0/xa2/XA1/a_1656_2090# 0 1.1f $ **FLOATING
C260 xbb0/xa2/XA1/a_1224_n110# 0 0.807f $ **FLOATING
C261 xbb0/xa2/XA1/a_792_2090# 0 1.1f $ **FLOATING
C262 xbb0/xa2/XA1/a_360_n110# 0 0.893f
C263 xbb0/xa2/XA1/a_n72_n110# 0 2.55f $ **FLOATING
C264 xbb0/xa2/N 0 3.45f
C265 xbb0/xa1/XA1/a_3816_n110# 0 2.55f
C266 xbb0/xa1/XA1/a_2952_n110# 0 0.893f $ **FLOATING
C267 xbb0/xa1/XA1/a_2520_2090# 0 1.1f $ **FLOATING
C268 xbb0/xa1/XA1/a_2088_n110# 0 0.807f $ **FLOATING
C269 xbb0/xa1/XA1/a_1656_2090# 0 1.1f $ **FLOATING
C270 xbb0/xa1/XA1/a_1224_n110# 0 0.807f $ **FLOATING
C271 xbb0/xa1/XA1/a_792_2090# 0 1.1f $ **FLOATING
C272 xbb0/xa1/XA1/a_360_n110# 0 0.893f
C273 xbb0/xa1/XA1/a_n72_n110# 0 2.55f $ **FLOATING
C274 xbb1/xa3/M8/a_324_334# 0 0.422f
C275 IBPSR_1U 0 17.1f
C276 xbb1/xa2/a_324_334# 0 0.358f
C277 xbb1/xa2/a_324_n18# 0 0.422f
.ends

