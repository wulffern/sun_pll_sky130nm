magic
tech sky130B
magscale 1 2
timestamp 1667257200
<< checkpaint >>
rect 0 0 4056 5936
<< locali >>
rect 3432 384 3672 5552
rect 384 384 3672 624
rect 384 5312 3672 5552
rect 384 384 624 5552
rect 3432 384 3672 5552
rect 3816 0 4056 5936
rect 0 0 4056 240
rect 0 5696 4056 5936
rect 0 0 240 5936
rect 3816 0 4056 5936
rect 1200 4786 1368 4846
rect 1368 4786 1428 4846
rect 2892 1706 3060 1766
rect 2892 1882 3060 1942
rect 3060 1706 3120 1942
rect 1170 914 1230 2734
rect 1632 4170 1800 4230
rect 1632 4346 1800 4406
rect 1800 4170 1860 4406
rect 1632 826 2004 886
rect 1632 2586 2004 2646
rect 2004 826 2064 2646
rect 1632 826 2004 886
rect 1632 4698 2004 4758
rect 2004 826 2064 4758
rect 2892 826 3264 886
rect 2892 1354 3264 1414
rect 3264 826 3324 1414
rect 2892 826 3264 886
rect 2892 2234 3264 2294
rect 3264 826 3324 2294
<< m1 >>
rect 1524 384 1740 886
rect 660 384 876 988
rect 2784 0 3000 886
rect 1920 0 2136 988
rect 2460 914 2628 974
rect 2628 1178 2892 1238
rect 1632 2410 2628 2470
rect 2460 1442 2628 1502
rect 2628 914 2688 2470
rect 2892 2058 3060 2118
rect 1632 4522 3060 4582
rect 2892 2410 3060 2470
rect 3060 2058 3120 4582
rect 1632 4874 1800 4934
rect 1800 4874 1860 4934
<< m2 >>
rect 0 1970 216 2030
rect 3840 4522 4056 4582
rect 0 4434 216 4494
rect 0 914 216 974
rect 3840 4874 4056 4934
rect 0 2322 216 2382
rect 0 4786 216 4846
rect 0 2322 216 2382
rect 2212 2292 2460 2368
rect 108 2322 2212 2398
rect 2212 2292 2288 2398
rect 0 4786 216 4846
rect 952 4786 1200 4862
rect 108 4786 952 4862
rect 952 4786 1028 4862
rect 0 914 216 974
rect 952 914 1200 990
rect 108 914 952 990
rect 952 914 1028 990
rect 3840 4522 4056 4582
rect 1632 4522 1804 4598
rect 1804 4522 3948 4598
rect 1804 4522 1880 4598
rect 3840 4874 4056 4934
rect 1632 4874 1804 4950
rect 1804 4874 3948 4950
rect 1804 4874 1880 4950
rect 0 1970 216 2030
rect 2212 1970 2460 2046
rect 108 1970 2212 2046
rect 2212 1970 2288 2046
rect 0 4434 216 4494
rect 952 4434 1200 4510
rect 108 4434 952 4510
rect 952 4434 1028 4510
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa1
transform 1 0 768 0 1 768
box 768 768 2028 2528
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM xa2
transform 1 0 768 0 1 2528
box 768 2528 2028 4288
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL xa3
transform 1 0 768 0 1 4288
box 768 4288 2028 4640
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA xa4
transform 1 0 768 0 1 4640
box 768 4640 2028 5168
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLCM xb1
transform -1 0 3288 0 1 768
box 3288 768 4548 1296
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLCM xb2
transform -1 0 3288 0 1 1296
box 3288 1296 4548 1824
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL xb3
transform -1 0 3288 0 1 1824
box 3288 1824 4548 2176
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL xb4
transform -1 0 3288 0 1 2176
box 3288 2176 4548 2528
use cut_M1M2_2x1 
transform 1 0 1540 0 1 826
box 1540 826 1724 894
use cut_M1M2_2x1 
transform 1 0 1540 0 1 384
box 1540 384 1724 452
use cut_M1M2_2x1 
transform 1 0 676 0 1 900
box 676 900 860 968
use cut_M1M2_2x1 
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M2_2x1 
transform 1 0 2800 0 1 826
box 2800 826 2984 894
use cut_M1M2_2x1 
transform 1 0 2800 0 1 0
box 2800 0 2984 68
use cut_M1M2_2x1 
transform 1 0 1936 0 1 900
box 1936 900 2120 968
use cut_M1M2_2x1 
transform 1 0 1936 0 1 0
box 1936 0 2120 68
use cut_M1M2_2x1 
transform 1 0 2352 0 1 914
box 2352 914 2536 982
use cut_M1M2_2x1 
transform 1 0 2784 0 1 1178
box 2784 1178 2968 1246
use cut_M1M2_2x1 
transform 1 0 1524 0 1 2410
box 1524 2410 1708 2478
use cut_M1M2_2x1 
transform 1 0 2352 0 1 1442
box 2352 1442 2536 1510
use cut_M1M2_2x1 
transform 1 0 2784 0 1 2058
box 2784 2058 2968 2126
use cut_M1M2_2x1 
transform 1 0 1524 0 1 4522
box 1524 4522 1708 4590
use cut_M1M2_2x1 
transform 1 0 2784 0 1 2410
box 2784 2410 2968 2478
use cut_M1M2_2x1 
transform 1 0 1524 0 1 4874
box 1524 4874 1708 4942
use cut_M1M3_2x1 
transform 1 0 2368 0 1 2284
box 2368 2284 2568 2360
use cut_M1M3_2x1 
transform 1 0 1108 0 1 4786
box 1108 4786 1308 4862
use cut_M1M3_2x1 
transform 1 0 1108 0 1 914
box 1108 914 1308 990
use cut_M1M3_2x1 
transform 1 0 1524 0 1 4522
box 1524 4522 1724 4598
use cut_M1M3_2x1 
transform 1 0 1524 0 1 4874
box 1524 4874 1724 4950
use cut_M1M3_2x1 
transform 1 0 2368 0 1 1970
box 2368 1970 2568 2046
use cut_M1M3_2x1 
transform 1 0 1108 0 1 4434
box 1108 4434 1308 4510
<< labels >>
flabel locali s 3432 384 3672 5552 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
flabel locali s 3816 0 4056 5936 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel m2 s 0 1970 216 2030 0 FreeSans 400 0 0 0 CP_UP_N
port 2 nsew
flabel m2 s 3840 4522 4056 4582 0 FreeSans 400 0 0 0 LPF
port 3 nsew
flabel m2 s 0 4434 216 4494 0 FreeSans 400 0 0 0 CP_DOWN
port 4 nsew
flabel m2 s 0 914 216 974 0 FreeSans 400 0 0 0 VBN
port 5 nsew
flabel m2 s 3840 4874 4056 4934 0 FreeSans 400 0 0 0 LPFZ
port 7 nsew
flabel m2 s 0 2322 216 2382 0 FreeSans 400 0 0 0 PWRUP_1V8
port 8 nsew
flabel m2 s 0 4786 216 4846 0 FreeSans 400 0 0 0 KICK
port 9 nsew
<< end >>
