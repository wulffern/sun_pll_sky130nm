magic
tech sky130B
magscale 1 1
timestamp 1720908000
<< checkpaint >>
rect 0 0 92 34
<< locali >>
rect 0 0 92 34
<< m1 >>
rect 0 0 92 34
<< viali >>
rect 6 3 86 31
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 92 34
<< end >>
