magic
tech sky130B
magscale 1 2
timestamp 1709161200
<< checkpaint >>
rect 0 0 6576 5408
<< locali >>
rect 5952 384 6192 5024
rect 384 384 6192 624
rect 384 4784 6192 5024
rect 384 384 624 5024
rect 5952 384 6192 5024
rect 6336 0 6576 5408
rect 0 0 6576 240
rect 0 5168 6576 5408
rect 0 0 240 5408
rect 6336 0 6576 5408
rect 4992 3526 5112 3586
rect 5112 3730 5376 3790
rect 5112 3526 5172 3790
rect 4944 3466 5052 3526
rect 4992 3878 5112 3938
rect 5112 4082 5376 4142
rect 5112 3878 5172 4142
rect 4944 3818 5052 3878
rect 4992 1766 5112 1826
rect 5112 1970 5376 2030
rect 5112 1766 5172 2030
rect 4944 1706 5052 1766
rect 4992 2118 5112 2178
rect 5112 2322 5376 2382
rect 5112 2118 5172 2382
rect 4944 2058 5052 2118
rect 4992 2470 5112 2530
rect 5112 2674 5376 2734
rect 5112 2470 5172 2734
rect 4944 2410 5052 2470
rect 4992 2822 5112 2882
rect 5112 3026 5376 3086
rect 5112 2822 5172 3086
rect 4944 2762 5052 2822
rect 4992 3174 5112 3234
rect 5112 3378 5376 3438
rect 5112 3174 5172 3438
rect 4944 3114 5052 3174
rect 4992 1414 5112 1474
rect 5112 1618 5376 1678
rect 5112 1414 5172 1678
rect 4944 1354 5052 1414
rect 1404 2118 1584 2178
rect 1200 2674 1404 2734
rect 1404 2118 1464 2734
rect 1524 2058 1632 2118
<< m3 >>
rect 1516 384 1732 2176
rect 5700 384 5916 988
rect 4844 384 5060 1472
rect 2308 0 2524 2176
rect 4060 4704 4260 5408
rect 4060 4704 4260 5408
rect 4052 768 4268 5408
<< m1 >>
rect 1404 1062 1584 1122
rect 1200 2322 1404 2382
rect 1404 1062 1464 2382
rect 1524 1002 1632 1062
rect 1524 5348 1740 5408
rect 5268 0 5484 60
rect 5268 0 5484 60
rect 5376 914 5544 974
rect 5376 0 5544 60
rect 5544 0 5604 974
rect 1524 5348 1740 5408
rect 1632 2762 1800 2822
rect 1632 5348 1800 5408
rect 1800 2762 1860 5408
<< m2 >>
rect 1200 1618 1372 1694
rect 1372 3466 4944 3542
rect 1372 1618 1448 3542
rect 952 914 1200 990
rect 952 3818 4944 3894
rect 952 914 1028 3894
rect 4944 4170 5116 4246
rect 5116 1266 5376 1342
rect 5116 1266 5192 4246
use SUN_PLL_LSCORE xa3 
transform 1 0 768 0 1 768
box 768 768 3288 2176
use SUNTR_IVX1_CV xa4 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 2176
box 768 2176 3288 2528
use SUNTR_IVX1_CV xa5 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 2528
box 768 2528 3288 2880
use SUNTR_TAPCELLB_CV xa6 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 2880
box 768 2880 3288 3232
use SUNTRB_NDX1_CV xb1 ../SUN_TRB_SKY130NM
transform -1 0 5808 0 1 768
box 5808 768 8328 1472
use SUNTRB_IVX1_CV xb2_0 ../SUN_TRB_SKY130NM
transform -1 0 5808 0 1 1472
box 5808 1472 8328 1824
use SUNTRB_IVX1_CV xb2_1 ../SUN_TRB_SKY130NM
transform -1 0 5808 0 1 1824
box 5808 1824 8328 2176
use SUNTRB_IVX1_CV xb2_2 ../SUN_TRB_SKY130NM
transform -1 0 5808 0 1 2176
box 5808 2176 8328 2528
use SUNTRB_IVX1_CV xb2_3 ../SUN_TRB_SKY130NM
transform -1 0 5808 0 1 2528
box 5808 2528 8328 2880
use SUNTRB_IVX1_CV xb2_4 ../SUN_TRB_SKY130NM
transform -1 0 5808 0 1 2880
box 5808 2880 8328 3232
use SUNTRB_IVX1_CV xb2_5 ../SUN_TRB_SKY130NM
transform -1 0 5808 0 1 3232
box 5808 3232 8328 3584
use SUNTRB_IVX1_CV xb2_6 ../SUN_TRB_SKY130NM
transform -1 0 5808 0 1 3584
box 5808 3584 8328 3936
use SUNTRB_IVX1_CV xb2_7 ../SUN_TRB_SKY130NM
transform -1 0 5808 0 1 3936
box 5808 3936 8328 4288
use SUNTRB_TAPCELLBAVSS_CV xb3 ../SUN_TRB_SKY130NM
transform -1 0 5808 0 1 4288
box 5808 4288 8328 4640
use cut_M1M4_2x1 xcut0 
transform 1 0 1524 0 1 384
box 1524 384 1724 460
use cut_M1M4_2x1 xcut1 
transform 1 0 5708 0 1 384
box 5708 384 5908 460
use cut_M1M4_2x1 xcut2 
transform 1 0 4852 0 1 384
box 4852 384 5052 460
use cut_M1M4_2x1 xcut3 
transform 1 0 2316 0 1 0
box 2316 0 2516 76
use cut_M1M2_2x1 xcut4 
transform 1 0 1556 0 1 1002
box 1556 1002 1740 1070
use cut_M1M2_2x1 xcut5 
transform 1 0 1124 0 1 2322
box 1124 2322 1308 2390
use cut_M1M3_2x1 xcut6 
transform 1 0 1092 0 1 1618
box 1092 1618 1292 1694
use cut_M1M3_2x1 xcut7 
transform 1 0 4836 0 1 3466
box 4836 3466 5036 3542
use cut_M1M3_2x1 xcut8 
transform 1 0 1108 0 1 914
box 1108 914 1308 990
use cut_M1M3_2x1 xcut9 
transform 1 0 4852 0 1 3818
box 4852 3818 5052 3894
use cut_M1M3_2x1 xcut10 
transform 1 0 4836 0 1 4170
box 4836 4170 5036 4246
use cut_M1M3_2x1 xcut11 
transform 1 0 5268 0 1 1266
box 5268 1266 5468 1342
use cut_M1M2_2x1 xcut12 
transform 1 0 5268 0 1 914
box 5268 914 5452 982
use cut_M1M2_2x1 xcut13 
transform 1 0 1524 0 1 2762
box 1524 2762 1708 2830
<< labels >>
flabel locali s 5952 384 6192 5024 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
flabel locali s 6336 0 6576 5408 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel m1 s 1524 5348 1740 5408 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel m3 s 4060 4704 4260 5408 0 FreeSans 400 0 0 0 VDD_ROSC
port 3 nsew signal bidirectional
flabel m1 s 5268 0 5484 60 0 FreeSans 400 0 0 0 PWRUP_1V8
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 6576 5408
<< end >>
