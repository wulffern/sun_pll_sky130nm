magic
tech sky130B
magscale 1 2
timestamp 1707433200
<< checkpaint >>
rect 0 0 4128 6640
<< locali >>
rect 3504 384 3744 6256
rect 384 384 3744 624
rect 384 6016 3744 6256
rect 384 384 624 6256
rect 3504 384 3744 6256
rect 3888 0 4128 6640
rect 0 0 4128 240
rect 0 6400 4128 6640
rect 0 0 240 6640
rect 3888 0 4128 6640
rect 1404 4758 1584 4818
rect 1200 5314 1404 5374
rect 1404 4758 1464 5374
rect 1524 4698 1632 4758
rect 1524 5226 1740 5286
rect 1524 5754 1740 5814
rect 1092 1266 1308 1326
rect 1524 1354 1740 1414
<< m1 >>
rect 1404 1766 1584 1826
rect 1200 1970 1404 2030
rect 1404 1766 1464 2030
rect 1524 1706 1632 1766
rect 1404 2118 1584 2178
rect 1200 2322 1404 2382
rect 1404 2118 1464 2382
rect 1524 2058 1632 2118
rect 1404 2470 1584 2530
rect 1404 2660 2604 2720
rect 1200 4258 1404 4318
rect 1404 2470 1464 4318
rect 1524 2410 1632 2470
rect 1404 4406 1584 4466
rect 1200 4610 1404 4670
rect 1404 4406 1464 4670
rect 1524 4346 1632 4406
rect 1200 5666 1368 5726
rect 1368 5226 1632 5286
rect 1368 5226 1428 5726
rect 972 1618 1200 1678
rect 972 1354 1632 1414
rect 972 4962 1200 5022
rect 972 1354 1032 5022
<< m3 >>
rect 1516 384 1732 5872
rect 1516 384 1732 3980
rect 2308 768 2524 6640
use SUNTR_TAPCELLB_CV xa1a ../SUN_TR_SKY130NM
transform 1 0 768 0 1 768
box 768 768 3288 1120
use SUNTR_IVX1_CV xa1b ../SUN_TR_SKY130NM
transform 1 0 768 0 1 1120
box 768 1120 3288 1472
use SUNTR_IVX1_CV xa1c ../SUN_TR_SKY130NM
transform 1 0 768 0 1 1472
box 768 1472 3288 1824
use SUNTR_IVX1_CV xa2 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 1824
box 768 1824 3288 2176
use SUNTR_IVX1_CV xa5a ../SUN_TR_SKY130NM
transform 1 0 768 0 1 2176
box 768 2176 3288 2528
use SUNTR_DCAPX1_CV xa5capb ../SUN_TR_SKY130NM
transform 1 0 768 0 1 2528
box 768 2528 3360 4112
use SUNTR_IVX1_CV xa6 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 4112
box 768 4112 3288 4464
use SUNTR_IVX1_CV xa7 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 4464
box 768 4464 3288 4816
use SUNTR_NRX1_CV xa8 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 4816
box 768 4816 3288 5520
use SUNTR_IVX1_CV xa9 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 5520
box 768 5520 3288 5872
use cut_M1M2_2x1 xcut0 
transform 1 0 1556 0 1 1706
box 1556 1706 1740 1774
use cut_M1M2_2x1 xcut1 
transform 1 0 1124 0 1 1970
box 1124 1970 1308 2038
use cut_M1M2_2x1 xcut2 
transform 1 0 1556 0 1 2058
box 1556 2058 1740 2126
use cut_M1M2_2x1 xcut3 
transform 1 0 1124 0 1 2322
box 1124 2322 1308 2390
use cut_M1M2_2x1 xcut4 
transform 1 0 1556 0 1 2410
box 1556 2410 1740 2478
use cut_M1M2_2x1 xcut5 
transform 1 0 2564 0 1 2660
box 2564 2660 2748 2728
use cut_M1M2_2x1 xcut6 
transform 1 0 1124 0 1 4258
box 1124 4258 1308 4326
use cut_M1M2_2x1 xcut7 
transform 1 0 1556 0 1 4346
box 1556 4346 1740 4414
use cut_M1M2_2x1 xcut8 
transform 1 0 1124 0 1 4610
box 1124 4610 1308 4678
use cut_M1M2_2x1 xcut9 
transform 1 0 1092 0 1 5666
box 1092 5666 1276 5734
use cut_M1M2_2x1 xcut10 
transform 1 0 1524 0 1 5226
box 1524 5226 1708 5294
use cut_M1M2_2x1 xcut11 
transform 1 0 1092 0 1 1618
box 1092 1618 1276 1686
use cut_M1M2_2x1 xcut12 
transform 1 0 1524 0 1 1354
box 1524 1354 1708 1422
use cut_M1M2_2x1 xcut13 
transform 1 0 1092 0 1 4962
box 1092 4962 1276 5030
use cut_M1M4_2x1 xcut14 
transform 1 0 1524 0 1 384
box 1524 384 1724 460
use cut_M1M4_2x1 xcut15 
transform 1 0 1524 0 1 3892
box 1524 3892 1724 3968
use cut_M1M4_2x1 xcut16 
transform 1 0 2316 0 1 6400
box 2316 6400 2516 6476
<< labels >>
flabel locali s 3504 384 3744 6256 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
flabel locali s 3888 0 4128 6640 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel locali s 1524 5226 1740 5286 0 FreeSans 400 0 0 0 KICK
port 2 nsew signal bidirectional
flabel locali s 1524 5754 1740 5814 0 FreeSans 400 0 0 0 KICK_N
port 3 nsew signal bidirectional
flabel locali s 1092 1266 1308 1326 0 FreeSans 400 0 0 0 PWRUP_1V8
port 4 nsew signal bidirectional
flabel locali s 1524 1354 1740 1414 0 FreeSans 400 0 0 0 PWRUP_1V8_N
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 4128 6640
<< end >>
