magic
tech sky130B
magscale 1 1
timestamp 1720908000
<< checkpaint >>
rect 0 0 100 38
<< locali >>
rect 0 0 92 34
<< m1 >>
rect 0 0 92 34
<< m2 >>
rect 0 0 100 38
<< viali >>
rect 6 3 86 31
<< v1 >>
rect 6 3 86 31
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 100 38
<< end >>
