magic
tech sky130B
magscale 1 1
timestamp 1720908000
<< checkpaint >>
rect 0 0 1260 704
<< locali >>
rect 813 117 843 235
rect 813 469 843 587
rect 828 645 912 675
rect 912 249 1044 279
rect 912 73 1044 103
rect 912 73 942 675
rect 432 469 516 499
rect 432 645 516 675
rect 516 469 546 675
rect 432 117 516 147
rect 432 293 516 323
rect 516 117 546 323
rect 216 73 300 103
rect 216 249 300 279
rect 300 73 330 279
rect 216 425 300 455
rect 216 601 300 631
rect 300 425 330 631
rect 432 293 516 323
rect 516 293 828 323
rect 516 293 546 323
rect 432 645 516 675
rect 516 645 828 675
rect 516 645 546 675
rect 378 645 486 675
rect 162 425 270 455
rect 162 73 270 103
rect 378 117 486 147
<< m1 >>
rect 828 293 912 323
rect 912 425 1044 455
rect 912 601 1044 631
rect 912 293 942 631
<< m3 >>
rect 774 0 874 704
rect 378 0 478 704
rect 774 0 874 704
rect 378 0 478 704
use SUNTR_NCHDL xb1_0 ../SUN_TR_SKY130NM
transform 1 0 0 0 1 0
box 0 0 630 176
use SUNTR_NCHDL xb1_1 ../SUN_TR_SKY130NM
transform 1 0 0 0 1 176
box 0 176 630 352
use SUNTR_NCHDL xb2_0 ../SUN_TR_SKY130NM
transform 1 0 0 0 1 352
box 0 352 630 528
use SUNTR_NCHDL xb2_1 ../SUN_TR_SKY130NM
transform 1 0 0 0 1 528
box 0 528 630 704
use SUNTR_PCHDL xc1a ../SUN_TR_SKY130NM
transform 1 0 630 0 1 0
box 630 0 1260 176
use SUNTR_PCHDL xc1b ../SUN_TR_SKY130NM
transform 1 0 630 0 1 176
box 630 176 1260 352
use SUNTR_PCHDL xc2a ../SUN_TR_SKY130NM
transform 1 0 630 0 1 352
box 630 352 1260 528
use SUNTR_PCHDL xc2b ../SUN_TR_SKY130NM
transform 1 0 630 0 1 528
box 630 528 1260 704
use cut_M1M2_2x1 xcut0 
transform 1 0 774 0 1 293
box 774 293 866 327
use cut_M1M2_2x1 xcut1 
transform 1 0 990 0 1 425
box 990 425 1082 459
use cut_M1M2_2x1 xcut2 
transform 1 0 990 0 1 601
box 990 601 1082 635
use cut_M1M4_2x1 xcut3 
transform 1 0 774 0 1 29
box 774 29 874 67
use cut_M1M4_2x1 xcut4 
transform 1 0 774 0 1 381
box 774 381 874 419
use cut_M1M4_2x1 xcut5 
transform 1 0 378 0 1 29
box 378 29 478 67
use cut_M1M4_2x1 xcut6 
transform 1 0 378 0 1 205
box 378 205 478 243
use cut_M1M4_2x1 xcut7 
transform 1 0 378 0 1 381
box 378 381 478 419
use cut_M1M4_2x1 xcut8 
transform 1 0 378 0 1 557
box 378 557 478 595
<< labels >>
flabel locali s 378 645 486 675 0 FreeSans 400 0 0 0 YN
port 3 nsew signal bidirectional
flabel locali s 162 425 270 455 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 162 73 270 103 0 FreeSans 400 0 0 0 AN
port 2 nsew signal bidirectional
flabel locali s 378 117 486 147 0 FreeSans 400 0 0 0 Y
port 4 nsew signal bidirectional
flabel m3 s 774 0 874 704 0 FreeSans 400 0 0 0 AVDD
port 5 nsew signal bidirectional
flabel m3 s 378 0 478 704 0 FreeSans 400 0 0 0 AVSS
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 704
<< end >>
