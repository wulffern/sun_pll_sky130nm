magic
tech sky130B
magscale 1 2
timestamp 1684706400
<< checkpaint >>
rect 0 0 200 76
<< locali >>
rect 0 0 184 68
<< m1 >>
rect 0 0 184 68
<< m2 >>
rect 0 0 200 76
<< viali >>
rect 12 6 172 62
<< v1 >>
rect 12 6 172 62
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 200 76
<< end >>
