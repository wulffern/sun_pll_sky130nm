magic
tech sky130B
magscale 1 2
timestamp 1680904800
<< checkpaint >>
rect 0 0 14712 11040
<< locali >>
rect 14088 384 14328 10656
rect 384 384 14328 624
rect 384 10416 14328 10656
rect 384 384 624 10656
rect 14088 384 14328 10656
rect 14472 0 14712 11040
rect 0 0 14712 240
rect 0 10800 14712 11040
rect 0 0 240 11040
rect 14472 0 14712 11040
rect 1632 2410 1800 2470
rect 1632 2586 1800 2646
rect 1632 3114 1800 3174
rect 1800 2410 1860 3174
rect 3252 826 3420 886
rect 3252 2410 3420 2470
rect 3252 3994 3420 4054
rect 3252 5578 3420 5638
rect 3252 7162 3420 7222
rect 3420 826 3480 7222
<< m1 >>
rect 1524 384 1740 886
rect 660 384 876 988
rect 660 384 876 2748
rect 660 384 876 3276
rect 3144 0 3360 886
rect 2280 0 2496 988
rect 2820 7250 2988 7310
rect 2988 1002 3252 1062
rect 2820 4082 2988 4142
rect 2820 5666 2988 5726
rect 1632 3290 2988 3350
rect 2988 1002 3048 7310
<< m3 >>
rect 8796 384 9012 812
rect 3252 4170 3432 4246
rect 3252 5754 3432 5830
rect 3252 7338 3432 7414
rect 3432 1604 8904 1680
rect 3432 2660 8904 2736
rect 3432 3716 8904 3792
rect 3432 4772 8904 4848
rect 3432 5828 8904 5904
rect 3432 6884 8904 6960
rect 3432 7940 8904 8016
rect 3432 8996 8904 9072
rect 3432 10052 8904 10128
rect 3432 1604 3508 10128
rect 8904 724 14196 800
rect 8904 1780 14196 1856
rect 8904 2836 14196 2912
rect 8904 3892 14196 3968
rect 8904 4948 14196 5024
rect 8904 6004 14196 6080
rect 8904 7060 14196 7136
rect 8904 8116 14196 8192
rect 8904 9172 14196 9248
rect 14196 724 14272 9248
<< m2 >>
rect 2820 914 2992 990
rect 1632 2762 2992 2838
rect 2992 2586 3252 2662
rect 2820 2498 2992 2574
rect 2992 914 3068 2838
rect 0 2674 216 2734
rect 0 3202 216 3262
rect 0 4170 216 4230
rect 0 914 216 974
rect 0 914 216 974
rect 952 914 1200 990
rect 108 914 952 990
rect 952 914 1028 990
rect 0 2674 216 2734
rect 952 2674 1200 2750
rect 108 2674 952 2750
rect 952 2674 1028 2750
rect 0 3202 216 3262
rect 952 3202 1200 3278
rect 108 3202 952 3278
rect 952 3202 1028 3278
rect 0 4170 216 4230
rect 3004 4170 3252 4246
rect 108 4170 3004 4246
rect 3004 4170 3080 4246
use ../SUN_TR_SKY130NM/SUNTR_NCHDLCM xa1
transform 1 0 768 0 1 768
box 768 768 2028 2528
use ../SUN_TR_SKY130NM/SUNTR_NCHDLA xa2
transform 1 0 768 0 1 2528
box 768 2528 2028 3056
use ../SUN_TR_SKY130NM/SUNTR_NCHDLA xa4
transform 1 0 768 0 1 3056
box 768 3056 2028 3584
use ../SUN_TR_SKY130NM/SUNTR_PCHDLA xc1
transform -1 0 3648 0 1 768
box 3648 768 4908 2352
use ../SUN_TR_SKY130NM/SUNTR_PCHDLA xc2
transform -1 0 3648 0 1 2352
box 3648 2352 4908 3936
use ../SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_0
transform -1 0 3648 0 1 3936
box 3648 3936 4908 5520
use ../SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_1
transform -1 0 3648 0 1 5520
box 3648 5520 4908 7104
use ../SUN_TR_SKY130NM/SUNTR_PCHDLA xc3_2
transform -1 0 3648 0 1 7104
box 3648 7104 4908 8688
use ../SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd2
transform 1 0 3792 0 1 768
box 3792 768 13944 1824
use ../SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd3_0
transform 1 0 3792 0 1 1824
box 3792 1824 13944 2880
use ../SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd3_1
transform 1 0 3792 0 1 2880
box 3792 2880 13944 3936
use ../SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd3_2
transform 1 0 3792 0 1 3936
box 3792 3936 13944 4992
use ../SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd3_3
transform 1 0 3792 0 1 4992
box 3792 4992 13944 6048
use ../SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd3_4
transform 1 0 3792 0 1 6048
box 3792 6048 13944 7104
use ../SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd3_5
transform 1 0 3792 0 1 7104
box 3792 7104 13944 8160
use ../SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd3_6
transform 1 0 3792 0 1 8160
box 3792 8160 13944 9216
use ../SUN_SAR9B_SKY130NM/SUNSAR_CAP_BSSW_CV xd3_7
transform 1 0 3792 0 1 9216
box 3792 9216 13944 10272
use cut_M1M2_2x1 xcut0
transform 1 0 1540 0 1 826
box 1540 826 1724 894
use cut_M1M2_2x1 xcut1
transform 1 0 1540 0 1 384
box 1540 384 1724 452
use cut_M1M2_2x1 xcut2
transform 1 0 676 0 1 900
box 676 900 860 968
use cut_M1M2_2x1 xcut3
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M2_2x1 xcut4
transform 1 0 676 0 1 2660
box 676 2660 860 2728
use cut_M1M2_2x1 xcut5
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M2_2x1 xcut6
transform 1 0 676 0 1 3188
box 676 3188 860 3256
use cut_M1M2_2x1 xcut7
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M4_2x1 xcut8
transform 1 0 8804 0 1 384
box 8804 384 9004 460
use cut_M1M2_2x1 xcut9
transform 1 0 3160 0 1 826
box 3160 826 3344 894
use cut_M1M2_2x1 xcut10
transform 1 0 3160 0 1 0
box 3160 0 3344 68
use cut_M1M2_2x1 xcut11
transform 1 0 2296 0 1 900
box 2296 900 2480 968
use cut_M1M2_2x1 xcut12
transform 1 0 2296 0 1 0
box 2296 0 2480 68
use cut_M1M2_2x1 xcut13
transform 1 0 2712 0 1 7250
box 2712 7250 2896 7318
use cut_M1M2_2x1 xcut14
transform 1 0 3144 0 1 1002
box 3144 1002 3328 1070
use cut_M1M2_2x1 xcut15
transform 1 0 2712 0 1 4082
box 2712 4082 2896 4150
use cut_M1M2_2x1 xcut16
transform 1 0 2712 0 1 5666
box 2712 5666 2896 5734
use cut_M1M2_2x1 xcut17
transform 1 0 1524 0 1 3290
box 1524 3290 1708 3358
use cut_M1M3_2x1 xcut18
transform 1 0 2712 0 1 914
box 2712 914 2912 990
use cut_M1M3_2x1 xcut19
transform 1 0 1524 0 1 2762
box 1524 2762 1724 2838
use cut_M1M3_2x1 xcut20
transform 1 0 3144 0 1 2586
box 3144 2586 3344 2662
use cut_M1M3_2x1 xcut21
transform 1 0 2712 0 1 2498
box 2712 2498 2912 2574
use cut_M1M4_2x1 xcut22
transform 1 0 3144 0 1 4170
box 3144 4170 3344 4246
use cut_M1M4_2x1 xcut23
transform 1 0 3144 0 1 5754
box 3144 5754 3344 5830
use cut_M1M4_2x1 xcut24
transform 1 0 3144 0 1 7338
box 3144 7338 3344 7414
use cut_M1M3_2x1 xcut25
transform 1 0 1108 0 1 914
box 1108 914 1308 990
use cut_M1M3_2x1 xcut26
transform 1 0 1108 0 1 2674
box 1108 2674 1308 2750
use cut_M1M3_2x1 xcut27
transform 1 0 1108 0 1 3202
box 1108 3202 1308 3278
<< labels >>
flabel locali s 14088 384 14328 10656 0 FreeSans 400 0 0 0 AVSS
port 6 nsew signal bidirectional
flabel locali s 14472 0 14712 11040 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel m2 s 0 2674 216 2734 0 FreeSans 400 0 0 0 VFB
port 2 nsew signal bidirectional
flabel m2 s 0 3202 216 3262 0 FreeSans 400 0 0 0 VI
port 3 nsew signal bidirectional
flabel m2 s 0 4170 216 4230 0 FreeSans 400 0 0 0 VO
port 4 nsew signal bidirectional
flabel m2 s 0 914 216 974 0 FreeSans 400 0 0 0 VBN
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 14712 11040
<< end >>
