magic
tech sky130B
timestamp 1681076574
<< locali >>
rect 0 5400 7356 5520
rect 0 120 120 5400
rect 192 5208 7164 5328
rect 192 312 312 5208
rect 1626 3581 1740 3611
rect 1710 2819 1740 3581
rect 1626 2789 1740 2819
rect 1710 2027 1740 2789
rect 1626 1997 1740 2027
rect 816 1557 930 1587
rect 900 1323 930 1557
rect 816 1293 930 1323
rect 900 1235 930 1293
rect 1710 1235 1740 1997
rect 816 1205 930 1235
rect 1626 1205 1740 1235
rect 1710 443 1740 1205
rect 1626 413 1740 443
rect 7044 312 7164 5208
rect 192 192 7164 312
rect 7236 120 7356 5400
rect 0 0 7356 120
<< metal1 >>
rect 1410 3625 1524 3655
rect 1494 2863 1524 3625
rect 1410 2833 1524 2863
rect 1494 2071 1524 2833
rect 1410 2041 1524 2071
rect 1494 1675 1524 2041
rect 816 1645 1524 1675
rect 330 192 438 1638
rect 1494 531 1524 1645
rect 1494 501 1626 531
rect 762 192 870 443
rect 1140 0 1248 494
rect 1572 0 1680 443
<< metal2 >>
rect 54 2115 1626 2123
rect 0 2085 1626 2115
rect 54 1631 600 1639
rect 0 1601 600 1631
rect 816 1381 1534 1419
rect 54 1367 600 1375
rect 0 1337 600 1367
rect 1496 1331 1534 1381
rect 1496 1293 1626 1331
rect 1496 1287 1534 1293
rect 1410 1249 1534 1287
rect 1496 495 1534 1249
rect 54 487 600 495
rect 0 457 600 487
rect 1410 457 1534 495
<< metal3 >>
rect 1716 5026 4452 5064
rect 1716 4536 1754 5026
rect 4452 4586 7136 4624
rect 1716 4498 4452 4536
rect 1716 4008 1754 4498
rect 7098 4096 7136 4586
rect 4452 4058 7136 4096
rect 1716 3970 4452 4008
rect 1716 3707 1754 3970
rect 1626 3669 1754 3707
rect 1716 3480 1754 3669
rect 7098 3568 7136 4058
rect 4452 3530 7136 3568
rect 1716 3442 4452 3480
rect 1716 2952 1754 3442
rect 7098 3040 7136 3530
rect 4452 3002 7136 3040
rect 1716 2915 4452 2952
rect 1626 2914 4452 2915
rect 1626 2877 1754 2914
rect 1716 2424 1754 2877
rect 7098 2512 7136 3002
rect 4452 2474 7136 2512
rect 1716 2386 4452 2424
rect 1716 2123 1754 2386
rect 1626 2085 1754 2123
rect 1716 1896 1754 2085
rect 7098 1984 7136 2474
rect 4452 1946 7136 1984
rect 1716 1858 4452 1896
rect 1716 1368 1754 1858
rect 7098 1456 7136 1946
rect 4452 1418 7136 1456
rect 1716 1330 4452 1368
rect 1716 840 1754 1330
rect 7098 928 7136 1418
rect 4452 890 7136 928
rect 1716 802 4452 840
rect 4398 400 4506 406
rect 7098 400 7136 890
rect 4398 362 7136 400
rect 4398 192 4506 362
use SUNTR_NCHDLCM  xa1 ../SUN_TR_SKY130NM
timestamp 1681076574
transform 1 0 384 0 1 384
box -90 -66 630 946
use SUNTR_NCHDLA  xa2 ../SUN_TR_SKY130NM
timestamp 1681076574
transform 1 0 384 0 1 1264
box -90 -66 630 330
use SUNTR_NCHDLA  xa4
timestamp 1681076574
transform 1 0 384 0 1 1528
box -90 -66 630 330
use SUNTR_PCHDLA  xc1 ../SUN_TR_SKY130NM
timestamp 1681076574
transform -1 0 1824 0 1 384
box 0 -66 720 858
use SUNTR_PCHDLA  xc2
timestamp 1681076574
transform -1 0 1824 0 1 1176
box 0 -66 720 858
use SUNTR_PCHDLA  xc3_0
timestamp 1681076574
transform -1 0 1824 0 1 1968
box 0 -66 720 858
use SUNTR_PCHDLA  xc3_1
timestamp 1681076574
transform -1 0 1824 0 1 2760
box 0 -66 720 858
use SUNTR_PCHDLA  xc3_2
timestamp 1681076574
transform -1 0 1824 0 1 3552
box 0 -66 720 858
use cut_M1M2_2x1  xcut0
timestamp 1680991200
transform 1 0 770 0 1 413
box 0 0 92 34
use cut_M1M2_2x1  xcut1
timestamp 1680991200
transform 1 0 770 0 1 192
box 0 0 92 34
use cut_M1M2_2x1  xcut2
timestamp 1680991200
transform 1 0 338 0 1 450
box 0 0 92 34
use cut_M1M2_2x1  xcut3
timestamp 1680991200
transform 1 0 338 0 1 192
box 0 0 92 34
use cut_M1M2_2x1  xcut4
timestamp 1680991200
transform 1 0 338 0 1 1330
box 0 0 92 34
use cut_M1M2_2x1  xcut5
timestamp 1680991200
transform 1 0 338 0 1 192
box 0 0 92 34
use cut_M1M2_2x1  xcut6
timestamp 1680991200
transform 1 0 338 0 1 1594
box 0 0 92 34
use cut_M1M2_2x1  xcut7
timestamp 1680991200
transform 1 0 338 0 1 192
box 0 0 92 34
use cut_M1M4_2x1  xcut8
timestamp 1680991200
transform 1 0 4402 0 1 192
box 0 0 100 38
use cut_M1M2_2x1  xcut9
timestamp 1680991200
transform 1 0 1580 0 1 413
box 0 0 92 34
use cut_M1M2_2x1  xcut10
timestamp 1680991200
transform 1 0 1580 0 1 0
box 0 0 92 34
use cut_M1M2_2x1  xcut11
timestamp 1680991200
transform 1 0 1148 0 1 450
box 0 0 92 34
use cut_M1M2_2x1  xcut12
timestamp 1680991200
transform 1 0 1148 0 1 0
box 0 0 92 34
use cut_M1M2_2x1  xcut13
timestamp 1680991200
transform 1 0 1356 0 1 3625
box 0 0 92 34
use cut_M1M2_2x1  xcut14
timestamp 1680991200
transform 1 0 1572 0 1 501
box 0 0 92 34
use cut_M1M2_2x1  xcut15
timestamp 1680991200
transform 1 0 1356 0 1 2041
box 0 0 92 34
use cut_M1M2_2x1  xcut16
timestamp 1680991200
transform 1 0 1356 0 1 2833
box 0 0 92 34
use cut_M1M2_2x1  xcut17
timestamp 1680991200
transform 1 0 762 0 1 1645
box 0 0 92 34
use cut_M1M3_2x1  xcut18
timestamp 1680991200
transform 1 0 1356 0 1 457
box 0 0 100 38
use cut_M1M3_2x1  xcut19
timestamp 1680991200
transform 1 0 762 0 1 1381
box 0 0 100 38
use cut_M1M3_2x1  xcut20
timestamp 1680991200
transform 1 0 1572 0 1 1293
box 0 0 100 38
use cut_M1M3_2x1  xcut21
timestamp 1680991200
transform 1 0 1356 0 1 1249
box 0 0 100 38
use cut_M1M4_2x1  xcut22
timestamp 1680991200
transform 1 0 1572 0 1 2085
box 0 0 100 38
use cut_M1M4_2x1  xcut23
timestamp 1680991200
transform 1 0 1572 0 1 2877
box 0 0 100 38
use cut_M1M4_2x1  xcut24
timestamp 1680991200
transform 1 0 1572 0 1 3669
box 0 0 100 38
use cut_M1M3_2x1  xcut25
timestamp 1680991200
transform 1 0 554 0 1 457
box 0 0 100 38
use cut_M1M3_2x1  xcut26
timestamp 1680991200
transform 1 0 554 0 1 1337
box 0 0 100 38
use cut_M1M3_2x1  xcut27
timestamp 1680991200
transform 1 0 554 0 1 1601
box 0 0 100 38
use SUNSAR_CAP_BSSW_CV  xd2 ../SUN_SAR9B_SKY130NM
timestamp 1680904800
transform 1 0 1896 0 1 384
box 54 -22 5058 462
use SUNSAR_CAP_BSSW_CV  xd3_0
timestamp 1680904800
transform 1 0 1896 0 1 912
box 54 -22 5058 462
use SUNSAR_CAP_BSSW_CV  xd3_1
timestamp 1680904800
transform 1 0 1896 0 1 1440
box 54 -22 5058 462
use SUNSAR_CAP_BSSW_CV  xd3_2
timestamp 1680904800
transform 1 0 1896 0 1 1968
box 54 -22 5058 462
use SUNSAR_CAP_BSSW_CV  xd3_3
timestamp 1680904800
transform 1 0 1896 0 1 2496
box 54 -22 5058 462
use SUNSAR_CAP_BSSW_CV  xd3_4
timestamp 1680904800
transform 1 0 1896 0 1 3024
box 54 -22 5058 462
use SUNSAR_CAP_BSSW_CV  xd3_5
timestamp 1680904800
transform 1 0 1896 0 1 3552
box 54 -22 5058 462
use SUNSAR_CAP_BSSW_CV  xd3_6
timestamp 1680904800
transform 1 0 1896 0 1 4080
box 54 -22 5058 462
use SUNSAR_CAP_BSSW_CV  xd3_7
timestamp 1680904800
transform 1 0 1896 0 1 4608
box 54 -22 5058 462
<< labels >>
flabel locali s 7044 192 7164 5328 0 FreeSans 200 0 0 0 AVSS
port 6 nsew signal bidirectional
flabel locali s 7236 0 7356 5520 0 FreeSans 200 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel metal2 s 0 1337 108 1367 0 FreeSans 200 0 0 0 VFB
port 2 nsew signal bidirectional
flabel metal2 s 0 1601 108 1631 0 FreeSans 200 0 0 0 VI
port 3 nsew signal bidirectional
flabel metal2 s 0 2085 108 2115 0 FreeSans 200 0 0 0 VO
port 4 nsew signal bidirectional
flabel metal2 s 0 457 108 487 0 FreeSans 200 0 0 0 VBN
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 7356 5520
<< end >>
