magic
tech sky130B
timestamp 1681076574
<< locali >>
rect 378 645 942 675
rect 216 601 330 631
rect 300 455 330 601
rect 516 499 546 645
rect 432 469 546 499
rect 813 469 843 587
rect 162 425 330 455
rect 432 293 828 323
rect 216 249 330 279
rect 300 103 330 249
rect 516 147 546 293
rect 912 279 942 645
rect 912 249 1044 279
rect 378 117 546 147
rect 813 117 843 235
rect 162 73 330 103
rect 912 103 942 249
rect 912 73 1044 103
<< metal1 >>
rect 912 601 1044 631
rect 912 455 942 601
rect 912 425 1044 455
rect 912 323 942 425
rect 828 293 942 323
<< metal3 >>
rect 378 0 478 704
rect 774 0 874 704
use SUNTR_NCHDL  xb1_0 ../SUN_TR_SKY130NM
timestamp 1680904800
transform 1 0 0 0 1 0
box -90 -66 630 242
use SUNTR_NCHDL  xb1_1
timestamp 1680904800
transform 1 0 0 0 1 176
box -90 -66 630 242
use SUNTR_NCHDL  xb2_0
timestamp 1680904800
transform 1 0 0 0 1 352
box -90 -66 630 242
use SUNTR_NCHDL  xb2_1
timestamp 1680904800
transform 1 0 0 0 1 528
box -90 -66 630 242
use SUNTR_PCHDL  xc1a ../SUN_TR_SKY130NM
timestamp 1680904800
transform 1 0 630 0 1 0
box 0 -66 720 242
use SUNTR_PCHDL  xc1b
timestamp 1680904800
transform 1 0 630 0 1 176
box 0 -66 720 242
use SUNTR_PCHDL  xc2a
timestamp 1680904800
transform 1 0 630 0 1 352
box 0 -66 720 242
use SUNTR_PCHDL  xc2b
timestamp 1680904800
transform 1 0 630 0 1 528
box 0 -66 720 242
use cut_M1M2_2x1  xcut0
timestamp 1680991200
transform 1 0 774 0 1 293
box 0 0 92 34
use cut_M1M2_2x1  xcut1
timestamp 1680991200
transform 1 0 990 0 1 425
box 0 0 92 34
use cut_M1M2_2x1  xcut2
timestamp 1680991200
transform 1 0 990 0 1 601
box 0 0 92 34
use cut_M1M4_2x1  xcut3
timestamp 1680991200
transform 1 0 774 0 1 29
box 0 0 100 38
use cut_M1M4_2x1  xcut4
timestamp 1680991200
transform 1 0 774 0 1 381
box 0 0 100 38
use cut_M1M4_2x1  xcut5
timestamp 1680991200
transform 1 0 378 0 1 29
box 0 0 100 38
use cut_M1M4_2x1  xcut6
timestamp 1680991200
transform 1 0 378 0 1 205
box 0 0 100 38
use cut_M1M4_2x1  xcut7
timestamp 1680991200
transform 1 0 378 0 1 381
box 0 0 100 38
use cut_M1M4_2x1  xcut8
timestamp 1680991200
transform 1 0 378 0 1 557
box 0 0 100 38
<< labels >>
flabel locali s 378 645 486 675 0 FreeSans 200 0 0 0 YN
port 3 nsew signal bidirectional
flabel locali s 162 425 270 455 0 FreeSans 200 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 162 73 270 103 0 FreeSans 200 0 0 0 AN
port 2 nsew signal bidirectional
flabel locali s 378 117 486 147 0 FreeSans 200 0 0 0 Y
port 4 nsew signal bidirectional
flabel metal3 s 774 0 874 704 0 FreeSans 200 0 0 0 AVDD
port 5 nsew signal bidirectional
flabel metal3 s 378 0 478 704 0 FreeSans 200 0 0 0 AVSS
port 6 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 704
<< end >>
