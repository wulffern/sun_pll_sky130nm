magic
tech sky130B
timestamp 1728046668
<< locali >>
rect 0 2584 3288 2704
rect 0 120 120 2584
rect 192 2392 3096 2512
rect 192 312 312 2392
rect 2556 2041 2688 2071
rect 2556 1969 2586 2041
rect 2496 1939 2586 1969
rect 2472 1909 2526 1939
rect 2556 1865 2688 1895
rect 2556 1793 2586 1865
rect 2496 1763 2586 1793
rect 2472 1733 2526 1763
rect 2556 1689 2688 1719
rect 2556 1617 2586 1689
rect 2496 1587 2586 1617
rect 2472 1557 2526 1587
rect 2556 1513 2688 1543
rect 2556 1441 2586 1513
rect 2496 1411 2586 1441
rect 2472 1381 2526 1411
rect 600 1337 732 1367
rect 702 1089 732 1337
rect 2556 1337 2688 1367
rect 2556 1265 2586 1337
rect 2496 1235 2586 1265
rect 2472 1205 2526 1235
rect 2556 1161 2688 1191
rect 2556 1089 2586 1161
rect 702 1059 792 1089
rect 2496 1059 2586 1089
rect 762 1029 816 1059
rect 2472 1029 2526 1059
rect 2556 985 2688 1015
rect 2556 913 2586 985
rect 2496 883 2586 913
rect 2472 853 2526 883
rect 2556 809 2688 839
rect 2556 737 2586 809
rect 2496 707 2586 737
rect 2472 677 2526 707
rect 2976 312 3096 2392
rect 192 192 3096 312
rect 3168 120 3288 2584
rect 0 0 3288 120
<< metal1 >>
rect 762 2674 930 2704
rect 900 1411 930 2674
rect 816 1381 930 1411
rect 600 1161 732 1191
rect 702 561 732 1161
rect 702 531 792 561
rect 762 501 816 531
rect 2688 457 2802 487
rect 2772 30 2802 457
rect 2634 0 2802 30
<< metal2 >>
rect 2472 2085 2596 2123
rect 476 1909 2472 1947
rect 476 495 514 1909
rect 686 1733 2472 1771
rect 686 847 724 1733
rect 600 809 724 847
rect 2558 671 2596 2085
rect 2558 633 2688 671
rect 476 457 600 495
<< metal3 >>
rect 758 192 866 1088
rect 1154 0 1262 1088
rect 2026 384 2134 2704
rect 2422 192 2530 736
rect 2850 192 2958 494
use SUN_PLL_LSCORE  xa3
timestamp 1728046668
transform 1 0 384 0 1 384
box -90 -66 1350 770
use SUNTR_IVX1_CV  xa4 ../SUN_TR_SKY130NM
timestamp 1728046668
transform 1 0 384 0 1 1088
box -90 -66 1350 242
use SUNTR_IVX1_CV  xa5
timestamp 1728046668
transform 1 0 384 0 1 1264
box -90 -66 1350 242
use SUNTR_TAPCELLB_CV  xa6 ../SUN_TR_SKY130NM
timestamp 1728046668
transform 1 0 384 0 1 1440
box -90 -66 1350 242
use SUNTRB_NDX1_CV  xb1 ../SUN_TRB_SKY130NM
timestamp 1728046668
transform -1 0 2904 0 1 384
box -90 -66 1350 418
use SUNTRB_IVX1_CV  xb2_0 ../SUN_TRB_SKY130NM
timestamp 1728046668
transform -1 0 2904 0 1 736
box -90 -66 1350 242
use SUNTRB_IVX1_CV  xb2_1
timestamp 1728046668
transform -1 0 2904 0 1 912
box -90 -66 1350 242
use SUNTRB_IVX1_CV  xb2_2
timestamp 1728046668
transform -1 0 2904 0 1 1088
box -90 -66 1350 242
use SUNTRB_IVX1_CV  xb2_3
timestamp 1728046668
transform -1 0 2904 0 1 1264
box -90 -66 1350 242
use SUNTRB_IVX1_CV  xb2_4
timestamp 1728046668
transform -1 0 2904 0 1 1440
box -90 -66 1350 242
use SUNTRB_IVX1_CV  xb2_5
timestamp 1728046668
transform -1 0 2904 0 1 1616
box -90 -66 1350 242
use SUNTRB_IVX1_CV  xb2_6
timestamp 1728046668
transform -1 0 2904 0 1 1792
box -90 -66 1350 242
use SUNTRB_IVX1_CV  xb2_7
timestamp 1728046668
transform -1 0 2904 0 1 1968
box -90 -66 1350 242
use SUNTRB_TAPCELLBAVSS_CV  xb3 ../SUN_TRB_SKY130NM
timestamp 1728046668
transform -1 0 2904 0 1 2144
box -90 -66 1350 242
use cut_M1M4_2x1  xcut0
timestamp 1720908000
transform 1 0 762 0 1 192
box 0 0 100 38
use cut_M1M4_2x1  xcut1
timestamp 1720908000
transform 1 0 2854 0 1 192
box 0 0 100 38
use cut_M1M4_2x1  xcut2
timestamp 1720908000
transform 1 0 2426 0 1 192
box 0 0 100 38
use cut_M1M4_2x1  xcut3
timestamp 1720908000
transform 1 0 1158 0 1 0
box 0 0 100 38
use cut_M1M2_2x1  xcut4
timestamp 1720908000
transform 1 0 778 0 1 501
box 0 0 92 34
use cut_M1M2_2x1  xcut5
timestamp 1720908000
transform 1 0 562 0 1 1161
box 0 0 92 34
use cut_M1M3_2x1  xcut6
timestamp 1720908000
transform 1 0 546 0 1 809
box 0 0 100 38
use cut_M1M3_2x1  xcut7
timestamp 1720908000
transform 1 0 2418 0 1 1733
box 0 0 100 38
use cut_M1M3_2x1  xcut8
timestamp 1720908000
transform 1 0 554 0 1 457
box 0 0 100 38
use cut_M1M3_2x1  xcut9
timestamp 1720908000
transform 1 0 2426 0 1 1909
box 0 0 100 38
use cut_M1M3_2x1  xcut10
timestamp 1720908000
transform 1 0 2418 0 1 2085
box 0 0 100 38
use cut_M1M3_2x1  xcut11
timestamp 1720908000
transform 1 0 2634 0 1 633
box 0 0 100 38
use cut_M1M2_2x1  xcut12
timestamp 1720908000
transform 1 0 2634 0 1 457
box 0 0 92 34
use cut_M1M2_2x1  xcut13
timestamp 1720908000
transform 1 0 762 0 1 1381
box 0 0 92 34
<< labels >>
flabel locali s 2976 192 3096 2512 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
flabel locali s 3168 0 3288 2704 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel metal1 s 762 2674 870 2704 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel metal3 s 2030 2352 2130 2704 0 FreeSans 400 0 0 0 VDD_ROSC
port 3 nsew signal bidirectional
flabel metal1 s 2634 0 2742 30 0 FreeSans 400 0 0 0 PWRUP_1V8
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 3288 2704
<< end >>
