*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/SUN_PLL_PFD_lpe.spi
#else
.include ../../../work/xsch/SUN_PLL_PFD.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

.param REF_PERIOD = 1/16e6
.param REF_HIGH = REF_PERIOD/2



.param FB_HIGH = FB_PERIOD/2


*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  AVSS  0     dc 0
VDD  AVDD 0  pwl 0 0 10n {AVDD}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

VREF CK_REF 0 dc 0 pulse (0 {AVDD} 0 {TRF} {TRF} {REF_HIGH} {REf_PERIOD})
VFB CK_FB 0 dc 0 pulse (0 {AVDD} 0 {TRF} {TRF} {FB_HIGH} {FB_PERIOD})


*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save CK_REF CK_FB CK_UP_N CP_DOWN v(xdut.cp_dup_n) v(xdut.cp_down_n) v(xdut.cp_up) v(xdut.cfb)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 10n 200n
write
quit


.endc

.end
