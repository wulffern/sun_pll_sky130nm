magic
tech sky130B
magscale 1 2
timestamp 1679854420
<< locali >>
rect -2000 66000 39000 67000
rect 2080 64696 2320 66000
rect 3680 64672 3920 66000
rect 5640 64000 5740 64120
rect -1980 63874 -1760 63880
rect -1980 63766 -1974 63874
rect -1866 63766 -1760 63874
rect -1980 63760 -1760 63766
rect 1816 57480 2056 59120
rect 5680 55014 6120 55020
rect 5680 54786 5686 55014
rect 5914 54786 6120 55014
rect 5680 54780 6120 54786
rect 5388 53780 5680 54020
rect 5388 51000 5628 51520
rect -2000 50414 39000 51000
rect -2000 50186 1386 50414
rect 1614 50186 39000 50414
rect -2000 50000 39000 50186
<< viali >>
rect 5520 64000 5640 64120
rect -1974 63766 -1866 63874
rect 5686 54786 5914 55014
rect 5680 53780 5920 54020
rect 1380 52384 1620 52624
rect 1386 50186 1614 50414
<< metal1 >>
rect 5520 65420 5640 65426
rect -1986 65300 -1980 65420
rect -1860 65300 -1854 65420
rect -1980 63874 -1860 65300
rect 5520 64126 5640 65300
rect 5508 64120 5652 64126
rect 5508 64000 5520 64120
rect 5640 64000 5652 64120
rect 5508 63994 5652 64000
rect -1980 63766 -1974 63874
rect -1866 63766 -1860 63874
rect -1980 63754 -1860 63766
rect -1996 59914 -1990 59974
rect -1930 59914 -1924 59974
rect -1990 58810 -1930 59914
rect -1990 58744 -1930 58750
rect 5680 55014 5920 55026
rect 5680 54786 5686 55014
rect 5914 54786 5920 55014
rect 5680 54032 5920 54786
rect 5674 54020 5926 54032
rect 5674 53780 5680 54020
rect 5920 53780 5926 54020
rect 5674 53768 5926 53780
rect 1368 52624 1632 52630
rect 1368 52384 1380 52624
rect 1620 52384 1632 52624
rect 1368 52378 1632 52384
rect 1380 50414 1620 52378
rect 1380 50186 1386 50414
rect 1614 50186 1620 50414
rect 1380 50174 1620 50186
<< via1 >>
rect -1980 65300 -1860 65420
rect 5520 65300 5640 65420
rect -1990 59914 -1930 59974
rect -1990 58750 -1930 58810
<< metal2 >>
rect -1980 65420 -1860 65426
rect -1860 65300 5520 65420
rect 5640 65300 5646 65420
rect -1980 65294 -1860 65300
rect -1957 63432 -1948 63488
rect -1892 63432 -1883 63488
rect -2100 61028 -1730 61030
rect -2107 60972 -2098 61028
rect -2042 60972 -1730 61028
rect -2100 60970 -1730 60972
rect -1990 59974 -1930 59980
rect -1990 59908 -1930 59914
rect -1996 58750 -1990 58810
rect -1930 58750 3790 58810
rect 2392 58230 2448 58237
rect -2109 58170 -2100 58230
rect -2040 58228 2450 58230
rect -2040 58172 2392 58228
rect 2448 58172 2450 58228
rect -2040 58170 2450 58172
rect 2392 58163 2448 58170
rect -1959 58030 -1950 58090
rect -1890 58088 2230 58090
rect -1890 58032 2172 58088
rect 2228 58032 2237 58088
rect -1890 58030 2230 58032
rect 1996 56874 2170 56934
rect 2230 56874 2239 56934
rect 1996 54762 2390 54822
rect 2450 54762 2459 54822
<< via2 >>
rect -1948 63432 -1892 63488
rect -2098 60972 -2042 61028
rect -2100 58170 -2040 58230
rect 2392 58172 2448 58228
rect -1950 58030 -1890 58090
rect 2172 58032 2228 58088
rect 2170 56874 2230 56934
rect 2390 54762 2450 54822
<< metal3 >>
rect -1953 63488 -1887 63493
rect -1953 63432 -1948 63488
rect -1892 63432 -1887 63488
rect -1953 63427 -1887 63432
rect -2103 61028 -2037 61033
rect -2103 60972 -2098 61028
rect -2042 60972 -2037 61028
rect -2103 60967 -2037 60972
rect -2100 58235 -2040 60967
rect -2105 58230 -2035 58235
rect -2105 58170 -2100 58230
rect -2040 58170 -2035 58230
rect -2105 58165 -2035 58170
rect -1950 58095 -1890 63427
rect 2387 58228 2453 58233
rect 2387 58172 2392 58228
rect 2448 58172 2453 58228
rect 2387 58167 2453 58172
rect -1955 58090 -1885 58095
rect -1955 58030 -1950 58090
rect -1890 58030 -1885 58090
rect -1955 58025 -1885 58030
rect 2167 58088 2233 58093
rect 2167 58032 2172 58088
rect 2228 58032 2233 58088
rect 2167 58027 2233 58032
rect 2170 56939 2230 58027
rect 2165 56934 2235 56939
rect 2165 56874 2170 56934
rect 2230 56874 2235 56934
rect 2165 56869 2235 56874
rect 2390 54827 2450 58167
rect 2385 54822 2455 54827
rect 2385 54762 2390 54822
rect 2450 54762 2455 54822
rect 2385 54757 2455 54762
use SUN_PLL_PFD  xaa0
timestamp 1679853665
transform 1 0 -2000 0 1 52000
box 0 0 4056 5760
use SUN_PLL_CP  xaa1
timestamp 1679853665
transform 1 0 -2000 0 1 59000
box 0 0 4344 5936
use SUN_PLL_KICK  xaa3
timestamp 1679854420
transform 1 0 3600 0 1 54400
box 0 0 4128 10512
use SUN_PLL_BUF  xaa4
timestamp 1679853665
transform 1 0 9000 0 1 52000
box 0 0 14712 11040
use SUN_PLL_ROSC  xaa5
timestamp 1679853665
transform 1 0 25000 0 1 60000
box 0 0 6576 5408
use SUN_PLL_DIVN  xaa6
timestamp 1679853665
transform 1 0 25000 0 1 52000
box 0 0 14136 7036
use SUN_PLL_LPF  xbb0
timestamp 1679853665
transform 1 0 -2000 0 1 69000
box 0 0 40552 49848
use SUN_PLL_BIAS  xbb1
timestamp 1679853665
transform 1 0 3600 0 1 51200
box 0 0 2028 2880
<< end >>
