magic
tech sky130B
magscale 1 2
timestamp 1684706400
<< checkpaint >>
rect 0 0 14784 13184
<< locali >>
rect 14160 384 14400 12768
rect 384 384 14400 624
rect 384 12528 14400 12768
rect 384 384 624 12768
rect 14160 384 14400 12768
rect 14544 0 14784 13152
rect 0 0 14784 240
rect 0 12912 14784 13152
rect 0 0 240 13152
rect 14544 0 14784 13152
rect 1632 2410 1800 2470
rect 1632 2586 1800 2646
rect 1632 4346 1800 4406
rect 1632 6106 1800 6166
rect 1632 7866 1800 7926
rect 1800 2410 1860 7926
rect 1170 6194 1230 8014
rect 1170 2674 1230 4494
rect 3324 914 3492 974
rect 3324 1442 3492 1502
rect 3324 1970 3492 2030
rect 3324 2498 3492 2558
rect 3324 3026 3492 3086
rect 3324 3554 3492 3614
rect 3324 4082 3492 4142
rect 3324 4610 3492 4670
rect 3324 5138 3492 5198
rect 3324 5666 3492 5726
rect 3324 6194 3492 6254
rect 3324 6722 3492 6782
rect 3324 7250 3492 7310
rect 3324 7778 3492 7838
rect 3324 8306 3492 8366
rect 3324 8834 3492 8894
rect 3324 9362 3492 9422
rect 3324 9890 3492 9950
rect 3324 10418 3492 10478
rect 3324 10946 3492 11006
rect 3324 11474 3492 11534
rect 3492 914 3552 11534
<< m1 >>
rect 1524 384 1740 886
rect 660 384 876 988
rect 3216 0 3432 974
rect 2352 0 2568 1076
rect 2892 11562 3060 11622
rect 1632 9450 3060 9510
rect 3060 3202 3324 3262
rect 3060 3730 3324 3790
rect 3060 4258 3324 4318
rect 3060 4786 3324 4846
rect 2892 5226 3060 5286
rect 2892 5754 3060 5814
rect 2892 6282 3060 6342
rect 2892 6810 3060 6870
rect 2892 7338 3060 7398
rect 2892 7866 3060 7926
rect 2892 8394 3060 8454
rect 2892 8922 3060 8982
rect 2892 9450 3060 9510
rect 2892 9978 3060 10038
rect 2892 10506 3060 10566
rect 2892 11034 3060 11094
rect 1632 7690 3060 7750
rect 3060 3202 3120 11622
rect 0 6194 216 6254
rect 0 6194 216 6254
rect 972 6194 1200 6254
rect 108 6194 972 6254
rect 972 6194 1032 6254
<< m3 >>
rect 8868 384 9084 812
rect 3324 5314 3504 5390
rect 3324 5842 3504 5918
rect 3324 6370 3504 6446
rect 3324 6898 3504 6974
rect 3324 7426 3504 7502
rect 3324 7954 3504 8030
rect 3324 8482 3504 8558
rect 3324 9010 3504 9086
rect 3324 9538 3504 9614
rect 3324 10066 3504 10142
rect 3324 10594 3504 10670
rect 3324 11122 3504 11198
rect 3324 11650 3504 11726
rect 3504 1604 8976 1680
rect 3504 2660 8976 2736
rect 3504 3716 8976 3792
rect 3504 4772 8976 4848
rect 3504 5828 8976 5904
rect 3504 6884 8976 6960
rect 3504 7940 8976 8016
rect 3504 8996 8976 9072
rect 3504 10052 8976 10128
rect 3504 11108 8976 11184
rect 3504 12164 8976 12240
rect 3504 1604 3580 12240
rect 8976 724 14268 800
rect 8976 1780 14268 1856
rect 8976 2836 14268 2912
rect 8976 3892 14268 3968
rect 8976 4948 14268 5024
rect 8976 6004 14268 6080
rect 8976 7060 14268 7136
rect 8976 8116 14268 8192
rect 8976 9172 14268 9248
rect 8976 10228 14268 10304
rect 8976 11284 14268 11360
rect 14268 724 14344 11360
rect 1092 13092 1308 13152
rect 3216 13108 3432 13168
rect 1092 13092 1308 13152
rect 944 2674 1200 2750
rect 944 13092 1200 13168
rect 944 2674 1020 13168
rect 3216 13108 3432 13168
rect 3324 5314 3504 5390
rect 3324 13108 3504 13184
rect 3504 5314 3580 13184
<< m2 >>
rect 2892 1002 3064 1078
rect 1632 5930 3064 6006
rect 3064 1090 3324 1166
rect 1632 4170 3064 4246
rect 3064 1618 3324 1694
rect 2892 1530 3064 1606
rect 3064 2146 3324 2222
rect 2892 2058 3064 2134
rect 3064 2674 3324 2750
rect 2892 2586 3064 2662
rect 2892 3114 3064 3190
rect 2892 3642 3064 3718
rect 2892 4170 3064 4246
rect 2892 4698 3064 4774
rect 3064 1002 3140 6006
rect 0 914 216 974
rect 0 914 216 974
rect 952 914 1200 990
rect 108 914 952 990
rect 952 914 1028 990
use SUNTR_NCHDLCM xa1 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 768
box 768 768 2028 2528
use SUNTR_NCHDLCM xa2_0 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 2528
box 768 2528 2028 4288
use SUNTR_NCHDLCM xa2_1 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 4288
box 768 4288 2028 6048
use SUNTR_NCHDLCM xa4_0 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 6048
box 768 6048 2028 7808
use SUNTR_NCHDLCM xa4_1 ../SUN_TR_SKY130NM
transform 1 0 768 0 1 7808
box 768 7808 2028 9568
use SUNTR_PCHL xc1_0 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 768
box 3720 768 4980 1296
use SUNTR_PCHL xc1_1 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 1296
box 3720 1296 4980 1824
use SUNTR_PCHL xc1_2 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 1824
box 3720 1824 4980 2352
use SUNTR_PCHL xc1_3 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 2352
box 3720 2352 4980 2880
use SUNTR_PCHL xc2_0 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 2880
box 3720 2880 4980 3408
use SUNTR_PCHL xc2_1 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 3408
box 3720 3408 4980 3936
use SUNTR_PCHL xc2_2 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 3936
box 3720 3936 4980 4464
use SUNTR_PCHL xc2_3 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 4464
box 3720 4464 4980 4992
use SUNTR_PCHL xc3_0 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 4992
box 3720 4992 4980 5520
use SUNTR_PCHL xc3_1 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 5520
box 3720 5520 4980 6048
use SUNTR_PCHL xc3_10 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 6048
box 3720 6048 4980 6576
use SUNTR_PCHL xc3_11 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 6576
box 3720 6576 4980 7104
use SUNTR_PCHL xc3_12 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 7104
box 3720 7104 4980 7632
use SUNTR_PCHL xc3_2 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 7632
box 3720 7632 4980 8160
use SUNTR_PCHL xc3_3 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 8160
box 3720 8160 4980 8688
use SUNTR_PCHL xc3_4 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 8688
box 3720 8688 4980 9216
use SUNTR_PCHL xc3_5 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 9216
box 3720 9216 4980 9744
use SUNTR_PCHL xc3_6 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 9744
box 3720 9744 4980 10272
use SUNTR_PCHL xc3_7 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 10272
box 3720 10272 4980 10800
use SUNTR_PCHL xc3_8 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 10800
box 3720 10800 4980 11328
use SUNTR_PCHL xc3_9 ../SUN_TR_SKY130NM
transform -1 0 3720 0 1 11328
box 3720 11328 4980 11856
use SUNSAR_CAP_BSSW_CV xd2 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 768
box 3864 768 14016 1824
use SUNSAR_CAP_BSSW_CV xd3_0 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 1824
box 3864 1824 14016 2880
use SUNSAR_CAP_BSSW_CV xd3_1 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 2880
box 3864 2880 14016 3936
use SUNSAR_CAP_BSSW_CV xd3_2 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 3936
box 3864 3936 14016 4992
use SUNSAR_CAP_BSSW_CV xd3_3 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 4992
box 3864 4992 14016 6048
use SUNSAR_CAP_BSSW_CV xd3_4 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 6048
box 3864 6048 14016 7104
use SUNSAR_CAP_BSSW_CV xd3_5 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 7104
box 3864 7104 14016 8160
use SUNSAR_CAP_BSSW_CV xd3_6 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 8160
box 3864 8160 14016 9216
use SUNSAR_CAP_BSSW_CV xd3_7 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 9216
box 3864 9216 14016 10272
use SUNSAR_CAP_BSSW_CV xd3_8 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 10272
box 3864 10272 14016 11328
use SUNSAR_CAP_BSSW_CV xd3_9 ../SUN_SAR9B_SKY130NM
transform 1 0 3864 0 1 11328
box 3864 11328 14016 12384
use cut_M1M2_2x1 xcut0 
transform 1 0 1540 0 1 826
box 1540 826 1724 894
use cut_M1M2_2x1 xcut1 
transform 1 0 1540 0 1 384
box 1540 384 1724 452
use cut_M1M2_2x1 xcut2 
transform 1 0 676 0 1 900
box 676 900 860 968
use cut_M1M2_2x1 xcut3 
transform 1 0 676 0 1 384
box 676 384 860 452
use cut_M1M4_2x1 xcut4 
transform 1 0 8876 0 1 384
box 8876 384 9076 460
use cut_M1M2_2x1 xcut5 
transform 1 0 3232 0 1 914
box 3232 914 3416 982
use cut_M1M2_2x1 xcut6 
transform 1 0 3232 0 1 0
box 3232 0 3416 68
use cut_M1M2_2x1 xcut7 
transform 1 0 2368 0 1 988
box 2368 988 2552 1056
use cut_M1M2_2x1 xcut8 
transform 1 0 2368 0 1 0
box 2368 0 2552 68
use cut_M1M2_2x1 xcut9 
transform 1 0 2784 0 1 11562
box 2784 11562 2968 11630
use cut_M1M2_2x1 xcut10 
transform 1 0 1524 0 1 9450
box 1524 9450 1708 9518
use cut_M1M2_2x1 xcut11 
transform 1 0 3216 0 1 3202
box 3216 3202 3400 3270
use cut_M1M2_2x1 xcut12 
transform 1 0 3216 0 1 3730
box 3216 3730 3400 3798
use cut_M1M2_2x1 xcut13 
transform 1 0 3216 0 1 4258
box 3216 4258 3400 4326
use cut_M1M2_2x1 xcut14 
transform 1 0 3216 0 1 4786
box 3216 4786 3400 4854
use cut_M1M2_2x1 xcut15 
transform 1 0 2784 0 1 5226
box 2784 5226 2968 5294
use cut_M1M2_2x1 xcut16 
transform 1 0 2784 0 1 5754
box 2784 5754 2968 5822
use cut_M1M2_2x1 xcut17 
transform 1 0 2784 0 1 6282
box 2784 6282 2968 6350
use cut_M1M2_2x1 xcut18 
transform 1 0 2784 0 1 6810
box 2784 6810 2968 6878
use cut_M1M2_2x1 xcut19 
transform 1 0 2784 0 1 7338
box 2784 7338 2968 7406
use cut_M1M2_2x1 xcut20 
transform 1 0 2784 0 1 7866
box 2784 7866 2968 7934
use cut_M1M2_2x1 xcut21 
transform 1 0 2784 0 1 8394
box 2784 8394 2968 8462
use cut_M1M2_2x1 xcut22 
transform 1 0 2784 0 1 8922
box 2784 8922 2968 8990
use cut_M1M2_2x1 xcut23 
transform 1 0 2784 0 1 9450
box 2784 9450 2968 9518
use cut_M1M2_2x1 xcut24 
transform 1 0 2784 0 1 9978
box 2784 9978 2968 10046
use cut_M1M2_2x1 xcut25 
transform 1 0 2784 0 1 10506
box 2784 10506 2968 10574
use cut_M1M2_2x1 xcut26 
transform 1 0 2784 0 1 11034
box 2784 11034 2968 11102
use cut_M1M2_2x1 xcut27 
transform 1 0 1524 0 1 7690
box 1524 7690 1708 7758
use cut_M1M3_2x1 xcut28 
transform 1 0 2784 0 1 1002
box 2784 1002 2984 1078
use cut_M1M3_2x1 xcut29 
transform 1 0 1524 0 1 5930
box 1524 5930 1724 6006
use cut_M1M3_2x1 xcut30 
transform 1 0 3216 0 1 1090
box 3216 1090 3416 1166
use cut_M1M3_2x1 xcut31 
transform 1 0 1524 0 1 4170
box 1524 4170 1724 4246
use cut_M1M3_2x1 xcut32 
transform 1 0 3216 0 1 1618
box 3216 1618 3416 1694
use cut_M1M3_2x1 xcut33 
transform 1 0 2784 0 1 1530
box 2784 1530 2984 1606
use cut_M1M3_2x1 xcut34 
transform 1 0 3216 0 1 2146
box 3216 2146 3416 2222
use cut_M1M3_2x1 xcut35 
transform 1 0 2784 0 1 2058
box 2784 2058 2984 2134
use cut_M1M3_2x1 xcut36 
transform 1 0 3216 0 1 2674
box 3216 2674 3416 2750
use cut_M1M3_2x1 xcut37 
transform 1 0 2784 0 1 2586
box 2784 2586 2984 2662
use cut_M1M3_2x1 xcut38 
transform 1 0 2784 0 1 3114
box 2784 3114 2984 3190
use cut_M1M3_2x1 xcut39 
transform 1 0 2784 0 1 3642
box 2784 3642 2984 3718
use cut_M1M3_2x1 xcut40 
transform 1 0 2784 0 1 4170
box 2784 4170 2984 4246
use cut_M1M3_2x1 xcut41 
transform 1 0 2784 0 1 4698
box 2784 4698 2984 4774
use cut_M1M4_2x1 xcut42 
transform 1 0 3216 0 1 5314
box 3216 5314 3416 5390
use cut_M1M4_2x1 xcut43 
transform 1 0 3216 0 1 5842
box 3216 5842 3416 5918
use cut_M1M4_2x1 xcut44 
transform 1 0 3216 0 1 6370
box 3216 6370 3416 6446
use cut_M1M4_2x1 xcut45 
transform 1 0 3216 0 1 6898
box 3216 6898 3416 6974
use cut_M1M4_2x1 xcut46 
transform 1 0 3216 0 1 7426
box 3216 7426 3416 7502
use cut_M1M4_2x1 xcut47 
transform 1 0 3216 0 1 7954
box 3216 7954 3416 8030
use cut_M1M4_2x1 xcut48 
transform 1 0 3216 0 1 8482
box 3216 8482 3416 8558
use cut_M1M4_2x1 xcut49 
transform 1 0 3216 0 1 9010
box 3216 9010 3416 9086
use cut_M1M4_2x1 xcut50 
transform 1 0 3216 0 1 9538
box 3216 9538 3416 9614
use cut_M1M4_2x1 xcut51 
transform 1 0 3216 0 1 10066
box 3216 10066 3416 10142
use cut_M1M4_2x1 xcut52 
transform 1 0 3216 0 1 10594
box 3216 10594 3416 10670
use cut_M1M4_2x1 xcut53 
transform 1 0 3216 0 1 11122
box 3216 11122 3416 11198
use cut_M1M4_2x1 xcut54 
transform 1 0 3216 0 1 11650
box 3216 11650 3416 11726
use cut_M1M3_2x1 xcut55 
transform 1 0 1108 0 1 914
box 1108 914 1308 990
use cut_M1M4_2x1 xcut56 
transform 1 0 1108 0 1 2674
box 1108 2674 1308 2750
use cut_M1M2_2x1 xcut57 
transform 1 0 1124 0 1 6194
box 1124 6194 1308 6262
<< labels >>
flabel locali s 14160 384 14400 12768 0 FreeSans 400 0 0 0 AVSS
port 6 nsew signal bidirectional
flabel locali s 14544 0 14784 13152 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel m3 s 1092 13092 1308 13152 0 FreeSans 400 0 0 0 VFB
port 2 nsew signal bidirectional
flabel m1 s 0 6194 216 6254 0 FreeSans 400 0 0 0 VI
port 3 nsew signal bidirectional
flabel m3 s 3216 13108 3432 13168 0 FreeSans 400 0 0 0 VO
port 4 nsew signal bidirectional
flabel m2 s 0 914 216 974 0 FreeSans 400 0 0 0 VBN
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 14784 13184
<< end >>
