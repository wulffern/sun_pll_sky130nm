* SUN_PLL_BUF

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/SUN_PLL_BUF_lpe.spi
.include ../../../work/lpe/SUN_PLL_BIAS_lpe.spi
#else
.include ../../../work/xsch/SUN_PLL_BIAS.spice
.include ../../../work/xsch/SUN_PLL_BUF.spice
#endif


*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
#ifdef Debug
.option reltol=1e-3 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-12
#else
*.option reltol=1e-5 srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-15
#endif

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  AVSS  0     dc 0
VDD  AVDD  AVSS  dc {AVDD}
VPWR PWRUP_1V8 AVSS dc {AVDD}
VCM VI 0 dc 1.2

IB 0 IBPSR_1U dc 1u

*-----------------------------------------------------------------
* Loop stability
*-----------------------------------------------------------------
.include ../../../../cpdk/ngspice/tian_subckt.lib
X999 LPI LPO loopgainprobe

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT0 IBPSR_1U AVSS AVSS SUN_PLL_BIAS
XDUT AVDD LPI VI LPO IBPSR_1U AVSS SUN_PLL_BUF

R1 LPO 0 100k
*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* SAVE
*----------------------------------------------------------------
.save V(X999.x) I(v.X999.Vi)
.save v(AVDD) v(VI) v(LPI) v(LPO) v(IBPSR_1U) v(AVSS)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit


optran 0 0 0 10n 1u 0
op
write {cicname}_op.raw

*----------------------------------------------------------------
* LSTB analysis
*----------------------------------------------------------------
* Set voltage AC to 1
ac dec 50 100 10G

* Set Current to 1
alter i.X999.Ii acmag=1
alter v.X999.Vi acmag=0
ac dec 50 100 10G

let lg_mag = db(tian_loop())
let lg_phase = 180*cph(tian_loop())/pi



write
quit
#endif

.endc

.end
