* SUN_PLL_BUF

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/SUN_PLL_BUF_lpe.spi
.include ../../../work/lpe/SUN_PLL_BIAS_lpe.spi
.include ../../../work/lpe/SUN_PLL_ROSC_lpe.spi
#else
.include ../../../work/xsch/SUN_PLL_BIAS.spice
.include ../../../work/xsch/SUN_PLL_BUF.spice
.include ../../../work/xsch/SUN_PLL_ROSC.spice
#endif


*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
#ifdef Debug
.option reltol=1e-3 srcsteps=1 ramptime=10n noopiter gmin=1e-12
#else
.option reltol=1e-3 srcsteps=1 ramptime=10n noopiter gmin=1e-15
#endif

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  AVSS  0  dc 0
VDD  AVDD  0  dc {AVDD}
VPWR PWRUP_1V8 0 dc {AVDD}
VI VI 0 pwl 0 {0} 6u {0} 20u {AVDD}

IB 0 IBPSR_1U dc 1u

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------

XDUT0 IBPSR_1U AVSS AVSS SUN_PLL_BIAS
XDUT AVDD VO VI VO IBPSR_1U AVSS SUN_PLL_BUF
XDUT2 AVDD CK VO PWRUP_1V8 AVSS SUN_PLL_ROSC


*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------

*----------------------------------------------------------------
* SAVE
*----------------------------------------------------------------
.save v(AVDD) v(VI) v(VO) v(IBPSR_1U) v(AVSS) v(XDUT.VGP) v(CK) i(vdd)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

tran 1n 20u
write
quit

.endc

.end


