

*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/SUN_PLL_lpe.spi
*.include ../../../work/lpe/SUN_PLL_BIAS_lpe.spi
*.include ../../../work/lpe/SUN_PLL_CP_lpe.spi
*.include ../../../work/lpe/SUN_PLL_DIVN_lpe.spi
*.include ../../../work/lpe/SUN_PLL_KICK_lpe.spi
*.include ../../../work/lpe/SUN_PLL_LPF_lpe.spi
*.include ../../../work/lpe/SUN_PLL_RCOSC_lpe.spi
*.include ../../../work/lpe/SUN_PLL_BUF_lpe.spi
*.include ../../../work/xsch/SUN_PLL.spice
#else
.include ../../../work/lpe/CAP_LPF_lpe.spi
.include ../../../work/lpe/SUNSAR_CAP_BSSW_CV_lpe.spi
.include ../../../work/xsch/SUN_PLL.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-15
#ifdef Debug
.option reltol=1e-3
#else
.option reltol=1e-4
#endif

.option TEMP=125
*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param PERIOD_CLK = 62.5n
.param PW_CLK = PERIOD_CLK/2

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  AVSS  0     dc 0
VDD  AVDD  AVSS  dc  {AVDD}
VPWR  PWRUP_1V8  AVSS pwl 0 0 1000n 0 1001n {AVDD}

IDC 0 IBPSR_1U  dc 1u


VCKREF CK_REF 0 dc 0 pulse (0 {AVDD} 0 {TRF} {TRF} {PW_CLK} {PERIOD_CLK})
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT AVDD AVSS PWRUP_1V8 CK_REF CK IBPSR_1U SUN_PLL

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* SAVE
*----------------------------------------------------------------

.save v(AVDD) v(AVSS) v(PWRUP_1V8) v(CK_REF) v(CK) v(IBPSR_1U)
.save v(XDUT.VDD_ROSC) v(XDUT.CP_UP_N) v(XDUT.CP_DOWN) v(XDUT.VLPF) v(XDUT.CK_FB) v(XDUT.KICK) v(XDUT.VLPFZ)
.save i(XDUT.AVDD) i(VDD)
.save v(XDUT.xaa3/KICK_N) v(XDUT.xaa3/KICK) v(XDUT.VLPZ)
.save v(XDUT.xaa4/VO)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=16
set color0=white
set color1=black
unset askquit

#ifdef Debug
tran 500p 3u
write
quit
#else
tran 200p 10u
write
quit
#endif

.endc

.end


