


*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option srcsteps=1 ramptime=10n noopiter keepopinfo gmin=1e-15
#ifdef Debug
.option reltol=1e-2
#else
.option reltol=1e-4
#endif


*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 100p

*.param PERIOD_CLK = 62.5n
.param PERIOD_CLK = 125n
.param PW_CLK = PERIOD_CLK/2

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  AVSS  0     dc 0
VDD  AVDD  AVSS  dc  {AVDD}
VPWR  PWRUP_1V8  AVSS pwl 0 0 1000n 0 1001n {AVDD}

IDC 0 IBPSR_1U  dc 1u


VCKREF CK_REF 0 dc 0 pulse (0 {AVDD} 0 {TRF} {TRF} {PW_CLK} {PERIOD_CLK})
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
*XDUT AVDD AVSS PWRUP_1V8 CK_REF CK IBPSR_1U SUN_PLL
.include ../xdut.spi

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* SAVE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save v(AVDD) v(AVSS) v(PWRUP_1V8) v(CK_REF) v(CK) v(IBPSR_1U)
.save v(XDUT.VDD_ROSC) v(XDUT.CP_UP_N) v(XDUT.CP_DOWN) v(XDUT.VLPF) v(XDUT.CK_FB) v(XDUT.KICK) v(XDUT.VLPFZ)
.save v(XDUT.*CP_DOWN) v(XDUT.*VLPF) v(XDUT.*CK_FB) v(XDUT.*KICK) v(XDUT.*VLPFZ)
.save i(XDUT.AVDD) i(VDD)
.save v(XDUT.xaa3/KICK_N) v(XDUT.xaa3/KICK) v(XDUT.VLPZ)
.save v(XDUT.xaa4/VO)
.save v(XDUT.xaa1/CP_UP_N) v(XDUT.xaa1/CP_DOWN)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=16
set color0=white
set color1=black
unset askquit

#ifdef Debug
tran 200p 3u
#else
tran 200p 15u
#endif
write
quit

rusage all

.endc

.end


