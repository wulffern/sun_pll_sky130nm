magic
tech sky130B
magscale 1 1
timestamp 1720908000
<< checkpaint >>
rect 0 0 100 38
<< m2 >>
rect 0 0 100 38
<< m3 >>
rect 0 0 100 38
<< v2 >>
rect 6 3 94 35
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 100 38
<< end >>
