magic
tech sky130B
magscale 1 2
timestamp 1680904800
<< checkpaint >>
rect 0 0 40552 49848
<< locali >>
rect 40252 0 40552 49848
rect 0 0 40552 300
rect 0 49548 40552 49848
rect 0 0 300 49848
rect 40252 0 40552 49848
rect 300 460 460 572
rect 300 5136 460 5248
rect 4516 8558 5092 8778
rect 1060 3882 1636 4102
<< m3 >>
rect 23120 0 23336 484
rect 39988 404 40328 480
rect 39988 1364 40328 1440
rect 39988 2324 40328 2400
rect 39988 3284 40328 3360
rect 39988 4244 40328 4320
rect 39988 5204 40328 5280
rect 39988 6164 40328 6240
rect 39988 7124 40328 7200
rect 39988 8084 40328 8160
rect 39988 9044 40328 9120
rect 39988 10004 40328 10080
rect 39988 10964 40328 11040
rect 39988 11924 40328 12000
rect 39988 12884 40328 12960
rect 39988 13844 40328 13920
rect 39988 14804 40328 14880
rect 39988 15764 40328 15840
rect 39988 16724 40328 16800
rect 39988 17684 40328 17760
rect 39988 18644 40328 18720
rect 39988 19604 40328 19680
rect 39988 20564 40328 20640
rect 39988 21524 40328 21600
rect 39988 22484 40328 22560
rect 39988 23444 40328 23520
rect 39988 24404 40328 24480
rect 39988 25364 40328 25440
rect 39988 26324 40328 26400
rect 39988 27284 40328 27360
rect 39988 28244 40328 28320
rect 39988 29204 40328 29280
rect 39988 30164 40328 30240
rect 39988 31124 40328 31200
rect 39988 32084 40328 32160
rect 39988 33044 40328 33120
rect 39988 34004 40328 34080
rect 39988 34964 40328 35040
rect 39988 35924 40328 36000
rect 39988 36884 40328 36960
rect 39988 37844 40328 37920
rect 39988 38804 40328 38880
rect 39988 39764 40328 39840
rect 39988 40724 40328 40800
rect 39988 41684 40328 41760
rect 39988 42644 40328 42720
rect 39988 43604 40328 43680
rect 39988 44564 40328 44640
rect 39988 45524 40328 45600
rect 39988 46484 40328 46560
rect 39988 47444 40328 47520
rect 39988 48404 40328 48480
<< m1 >>
rect 1152 8558 1508 8618
rect 1508 3882 4608 3942
rect 1508 3882 1568 8618
rect 4608 8558 4760 8618
rect 4760 4084 6568 4144
rect 4760 5044 6568 5104
rect 4760 6004 6568 6064
rect 4760 6964 6568 7024
rect 4760 7924 6568 7984
rect 4760 8884 6568 8944
rect 4760 9844 6568 9904
rect 4760 10804 6568 10864
rect 4760 11764 6568 11824
rect 4760 12724 6568 12784
rect 4760 13684 6568 13744
rect 4760 14644 6568 14704
rect 4760 15604 6568 15664
rect 4760 16564 6568 16624
rect 4760 17524 6568 17584
rect 4760 18484 6568 18544
rect 4760 19444 6568 19504
rect 4760 20404 6568 20464
rect 4760 21364 6568 21424
rect 4760 22324 6568 22384
rect 4760 23284 6568 23344
rect 4760 24244 6568 24304
rect 4760 25204 6568 25264
rect 4760 26164 6568 26224
rect 4760 27124 6568 27184
rect 4760 28084 6568 28144
rect 4760 29044 6568 29104
rect 4760 30004 6568 30064
rect 4760 30964 6568 31024
rect 4760 31924 6568 31984
rect 4760 32884 6568 32944
rect 4760 33844 6568 33904
rect 4760 34804 6568 34864
rect 4760 35764 6568 35824
rect 4760 36724 6568 36784
rect 4760 37684 6568 37744
rect 4760 38644 6568 38704
rect 4760 39604 6568 39664
rect 4760 40564 6568 40624
rect 4760 41524 6568 41584
rect 4760 42484 6568 42544
rect 4760 43444 6568 43504
rect 4760 44404 6568 44464
rect 4760 45364 6568 45424
rect 4760 46324 6568 46384
rect 4760 47284 6568 47344
rect 4760 48244 6568 48304
rect 4760 49204 6568 49264
rect 4760 4084 4820 49264
<< m2 >>
rect 1160 3882 1324 3958
rect 1324 1204 6568 1280
rect 1324 2164 6568 2240
rect 1324 3124 6568 3200
rect 1324 1204 1400 3958
use ../SUN_TR_SKY130NM/SUNTR_RPPO8 xa1
transform 1 0 444 0 1 444
box 444 444 5708 4680
use ../SUN_TR_SKY130NM/SUNTR_RPPO8 xa2
transform 1 0 444 0 1 5120
box 444 5120 5708 9356
use CAP_LPF xb1
transform -1 0 40108 0 1 444
box 40108 444 73788 1404
use CAP_LPF xb2_0
transform -1 0 40108 0 1 1404
box 40108 1404 73788 2364
use CAP_LPF xb2_1
transform -1 0 40108 0 1 2364
box 40108 2364 73788 3324
use CAP_LPF xb3_0
transform -1 0 40108 0 1 3324
box 40108 3324 73788 4284
use CAP_LPF xb3_1
transform -1 0 40108 0 1 4284
box 40108 4284 73788 5244
use CAP_LPF xb3_10
transform -1 0 40108 0 1 5244
box 40108 5244 73788 6204
use CAP_LPF xb3_11
transform -1 0 40108 0 1 6204
box 40108 6204 73788 7164
use CAP_LPF xb3_12
transform -1 0 40108 0 1 7164
box 40108 7164 73788 8124
use CAP_LPF xb3_13
transform -1 0 40108 0 1 8124
box 40108 8124 73788 9084
use CAP_LPF xb3_14
transform -1 0 40108 0 1 9084
box 40108 9084 73788 10044
use CAP_LPF xb3_15
transform -1 0 40108 0 1 10044
box 40108 10044 73788 11004
use CAP_LPF xb3_16
transform -1 0 40108 0 1 11004
box 40108 11004 73788 11964
use CAP_LPF xb3_17
transform -1 0 40108 0 1 11964
box 40108 11964 73788 12924
use CAP_LPF xb3_18
transform -1 0 40108 0 1 12924
box 40108 12924 73788 13884
use CAP_LPF xb3_19
transform -1 0 40108 0 1 13884
box 40108 13884 73788 14844
use CAP_LPF xb3_2
transform -1 0 40108 0 1 14844
box 40108 14844 73788 15804
use CAP_LPF xb3_20
transform -1 0 40108 0 1 15804
box 40108 15804 73788 16764
use CAP_LPF xb3_21
transform -1 0 40108 0 1 16764
box 40108 16764 73788 17724
use CAP_LPF xb3_22
transform -1 0 40108 0 1 17724
box 40108 17724 73788 18684
use CAP_LPF xb3_23
transform -1 0 40108 0 1 18684
box 40108 18684 73788 19644
use CAP_LPF xb3_24
transform -1 0 40108 0 1 19644
box 40108 19644 73788 20604
use CAP_LPF xb3_25
transform -1 0 40108 0 1 20604
box 40108 20604 73788 21564
use CAP_LPF xb3_26
transform -1 0 40108 0 1 21564
box 40108 21564 73788 22524
use CAP_LPF xb3_27
transform -1 0 40108 0 1 22524
box 40108 22524 73788 23484
use CAP_LPF xb3_28
transform -1 0 40108 0 1 23484
box 40108 23484 73788 24444
use CAP_LPF xb3_29
transform -1 0 40108 0 1 24444
box 40108 24444 73788 25404
use CAP_LPF xb3_3
transform -1 0 40108 0 1 25404
box 40108 25404 73788 26364
use CAP_LPF xb3_30
transform -1 0 40108 0 1 26364
box 40108 26364 73788 27324
use CAP_LPF xb3_31
transform -1 0 40108 0 1 27324
box 40108 27324 73788 28284
use CAP_LPF xb3_32
transform -1 0 40108 0 1 28284
box 40108 28284 73788 29244
use CAP_LPF xb3_33
transform -1 0 40108 0 1 29244
box 40108 29244 73788 30204
use CAP_LPF xb3_34
transform -1 0 40108 0 1 30204
box 40108 30204 73788 31164
use CAP_LPF xb3_35
transform -1 0 40108 0 1 31164
box 40108 31164 73788 32124
use CAP_LPF xb3_36
transform -1 0 40108 0 1 32124
box 40108 32124 73788 33084
use CAP_LPF xb3_37
transform -1 0 40108 0 1 33084
box 40108 33084 73788 34044
use CAP_LPF xb3_38
transform -1 0 40108 0 1 34044
box 40108 34044 73788 35004
use CAP_LPF xb3_39
transform -1 0 40108 0 1 35004
box 40108 35004 73788 35964
use CAP_LPF xb3_4
transform -1 0 40108 0 1 35964
box 40108 35964 73788 36924
use CAP_LPF xb3_40
transform -1 0 40108 0 1 36924
box 40108 36924 73788 37884
use CAP_LPF xb3_41
transform -1 0 40108 0 1 37884
box 40108 37884 73788 38844
use CAP_LPF xb3_42
transform -1 0 40108 0 1 38844
box 40108 38844 73788 39804
use CAP_LPF xb3_43
transform -1 0 40108 0 1 39804
box 40108 39804 73788 40764
use CAP_LPF xb3_44
transform -1 0 40108 0 1 40764
box 40108 40764 73788 41724
use CAP_LPF xb3_45
transform -1 0 40108 0 1 41724
box 40108 41724 73788 42684
use CAP_LPF xb3_46
transform -1 0 40108 0 1 42684
box 40108 42684 73788 43644
use CAP_LPF xb3_47
transform -1 0 40108 0 1 43644
box 40108 43644 73788 44604
use CAP_LPF xb3_5
transform -1 0 40108 0 1 44604
box 40108 44604 73788 45564
use CAP_LPF xb3_6
transform -1 0 40108 0 1 45564
box 40108 45564 73788 46524
use CAP_LPF xb3_7
transform -1 0 40108 0 1 46524
box 40108 46524 73788 47484
use CAP_LPF xb3_8
transform -1 0 40108 0 1 47484
box 40108 47484 73788 48444
use CAP_LPF xb3_9
transform -1 0 40108 0 1 48444
box 40108 48444 73788 49404
use cut_M1M4_2x1 xcut0
transform 1 0 23128 0 1 0
box 23128 0 23328 76
use cut_M1M2_2x1 xcut1
transform 1 0 1060 0 1 8558
box 1060 8558 1244 8626
use cut_M1M2_2x1 xcut2
transform 1 0 4516 0 1 3882
box 4516 3882 4700 3950
use cut_M1M2_2x1 xcut3
transform 1 0 4516 0 1 8558
box 4516 8558 4700 8626
use cut_M2M4_2x1 xcut4
transform 1 0 6468 0 1 4084
box 6468 4084 6668 4160
use cut_M2M4_2x1 xcut5
transform 1 0 6468 0 1 5044
box 6468 5044 6668 5120
use cut_M2M4_2x1 xcut6
transform 1 0 6468 0 1 6004
box 6468 6004 6668 6080
use cut_M2M4_2x1 xcut7
transform 1 0 6468 0 1 6964
box 6468 6964 6668 7040
use cut_M2M4_2x1 xcut8
transform 1 0 6468 0 1 7924
box 6468 7924 6668 8000
use cut_M2M4_2x1 xcut9
transform 1 0 6468 0 1 8884
box 6468 8884 6668 8960
use cut_M2M4_2x1 xcut10
transform 1 0 6468 0 1 9844
box 6468 9844 6668 9920
use cut_M2M4_2x1 xcut11
transform 1 0 6468 0 1 10804
box 6468 10804 6668 10880
use cut_M2M4_2x1 xcut12
transform 1 0 6468 0 1 11764
box 6468 11764 6668 11840
use cut_M2M4_2x1 xcut13
transform 1 0 6468 0 1 12724
box 6468 12724 6668 12800
use cut_M2M4_2x1 xcut14
transform 1 0 6468 0 1 13684
box 6468 13684 6668 13760
use cut_M2M4_2x1 xcut15
transform 1 0 6468 0 1 14644
box 6468 14644 6668 14720
use cut_M2M4_2x1 xcut16
transform 1 0 6468 0 1 15604
box 6468 15604 6668 15680
use cut_M2M4_2x1 xcut17
transform 1 0 6468 0 1 16564
box 6468 16564 6668 16640
use cut_M2M4_2x1 xcut18
transform 1 0 6468 0 1 17524
box 6468 17524 6668 17600
use cut_M2M4_2x1 xcut19
transform 1 0 6468 0 1 18484
box 6468 18484 6668 18560
use cut_M2M4_2x1 xcut20
transform 1 0 6468 0 1 19444
box 6468 19444 6668 19520
use cut_M2M4_2x1 xcut21
transform 1 0 6468 0 1 20404
box 6468 20404 6668 20480
use cut_M2M4_2x1 xcut22
transform 1 0 6468 0 1 21364
box 6468 21364 6668 21440
use cut_M2M4_2x1 xcut23
transform 1 0 6468 0 1 22324
box 6468 22324 6668 22400
use cut_M2M4_2x1 xcut24
transform 1 0 6468 0 1 23284
box 6468 23284 6668 23360
use cut_M2M4_2x1 xcut25
transform 1 0 6468 0 1 24244
box 6468 24244 6668 24320
use cut_M2M4_2x1 xcut26
transform 1 0 6468 0 1 25204
box 6468 25204 6668 25280
use cut_M2M4_2x1 xcut27
transform 1 0 6468 0 1 26164
box 6468 26164 6668 26240
use cut_M2M4_2x1 xcut28
transform 1 0 6468 0 1 27124
box 6468 27124 6668 27200
use cut_M2M4_2x1 xcut29
transform 1 0 6468 0 1 28084
box 6468 28084 6668 28160
use cut_M2M4_2x1 xcut30
transform 1 0 6468 0 1 29044
box 6468 29044 6668 29120
use cut_M2M4_2x1 xcut31
transform 1 0 6468 0 1 30004
box 6468 30004 6668 30080
use cut_M2M4_2x1 xcut32
transform 1 0 6468 0 1 30964
box 6468 30964 6668 31040
use cut_M2M4_2x1 xcut33
transform 1 0 6468 0 1 31924
box 6468 31924 6668 32000
use cut_M2M4_2x1 xcut34
transform 1 0 6468 0 1 32884
box 6468 32884 6668 32960
use cut_M2M4_2x1 xcut35
transform 1 0 6468 0 1 33844
box 6468 33844 6668 33920
use cut_M2M4_2x1 xcut36
transform 1 0 6468 0 1 34804
box 6468 34804 6668 34880
use cut_M2M4_2x1 xcut37
transform 1 0 6468 0 1 35764
box 6468 35764 6668 35840
use cut_M2M4_2x1 xcut38
transform 1 0 6468 0 1 36724
box 6468 36724 6668 36800
use cut_M2M4_2x1 xcut39
transform 1 0 6468 0 1 37684
box 6468 37684 6668 37760
use cut_M2M4_2x1 xcut40
transform 1 0 6468 0 1 38644
box 6468 38644 6668 38720
use cut_M2M4_2x1 xcut41
transform 1 0 6468 0 1 39604
box 6468 39604 6668 39680
use cut_M2M4_2x1 xcut42
transform 1 0 6468 0 1 40564
box 6468 40564 6668 40640
use cut_M2M4_2x1 xcut43
transform 1 0 6468 0 1 41524
box 6468 41524 6668 41600
use cut_M2M4_2x1 xcut44
transform 1 0 6468 0 1 42484
box 6468 42484 6668 42560
use cut_M2M4_2x1 xcut45
transform 1 0 6468 0 1 43444
box 6468 43444 6668 43520
use cut_M2M4_2x1 xcut46
transform 1 0 6468 0 1 44404
box 6468 44404 6668 44480
use cut_M2M4_2x1 xcut47
transform 1 0 6468 0 1 45364
box 6468 45364 6668 45440
use cut_M2M4_2x1 xcut48
transform 1 0 6468 0 1 46324
box 6468 46324 6668 46400
use cut_M2M4_2x1 xcut49
transform 1 0 6468 0 1 47284
box 6468 47284 6668 47360
use cut_M2M4_2x1 xcut50
transform 1 0 6468 0 1 48244
box 6468 48244 6668 48320
use cut_M2M4_2x1 xcut51
transform 1 0 6468 0 1 49204
box 6468 49204 6668 49280
use cut_M1M3_2x1 xcut52
transform 1 0 1060 0 1 3882
box 1060 3882 1260 3958
use cut_M3M4_2x1 xcut53
transform 1 0 6468 0 1 1204
box 6468 1204 6668 1280
use cut_M3M4_2x1 xcut54
transform 1 0 6468 0 1 2164
box 6468 2164 6668 2240
use cut_M3M4_2x1 xcut55
transform 1 0 6468 0 1 3124
box 6468 3124 6668 3200
use cut_M1M4_1x2 xcut56
transform 1 0 40252 0 1 0
box 40252 0 40328 200
use cut_M1M4_1x2 xcut57
transform 1 0 40252 0 1 404
box 40252 404 40328 604
use cut_M1M4_1x2 xcut58
transform 1 0 40252 0 1 1364
box 40252 1364 40328 1564
use cut_M1M4_1x2 xcut59
transform 1 0 40252 0 1 2324
box 40252 2324 40328 2524
use cut_M1M4_1x2 xcut60
transform 1 0 40252 0 1 3284
box 40252 3284 40328 3484
use cut_M1M4_1x2 xcut61
transform 1 0 40252 0 1 4244
box 40252 4244 40328 4444
use cut_M1M4_1x2 xcut62
transform 1 0 40252 0 1 5204
box 40252 5204 40328 5404
use cut_M1M4_1x2 xcut63
transform 1 0 40252 0 1 6164
box 40252 6164 40328 6364
use cut_M1M4_1x2 xcut64
transform 1 0 40252 0 1 7124
box 40252 7124 40328 7324
use cut_M1M4_1x2 xcut65
transform 1 0 40252 0 1 8084
box 40252 8084 40328 8284
use cut_M1M4_1x2 xcut66
transform 1 0 40252 0 1 9044
box 40252 9044 40328 9244
use cut_M1M4_1x2 xcut67
transform 1 0 40252 0 1 10004
box 40252 10004 40328 10204
use cut_M1M4_1x2 xcut68
transform 1 0 40252 0 1 10964
box 40252 10964 40328 11164
use cut_M1M4_1x2 xcut69
transform 1 0 40252 0 1 11924
box 40252 11924 40328 12124
use cut_M1M4_1x2 xcut70
transform 1 0 40252 0 1 12884
box 40252 12884 40328 13084
use cut_M1M4_1x2 xcut71
transform 1 0 40252 0 1 13844
box 40252 13844 40328 14044
use cut_M1M4_1x2 xcut72
transform 1 0 40252 0 1 14804
box 40252 14804 40328 15004
use cut_M1M4_1x2 xcut73
transform 1 0 40252 0 1 15764
box 40252 15764 40328 15964
use cut_M1M4_1x2 xcut74
transform 1 0 40252 0 1 16724
box 40252 16724 40328 16924
use cut_M1M4_1x2 xcut75
transform 1 0 40252 0 1 17684
box 40252 17684 40328 17884
use cut_M1M4_1x2 xcut76
transform 1 0 40252 0 1 18644
box 40252 18644 40328 18844
use cut_M1M4_1x2 xcut77
transform 1 0 40252 0 1 19604
box 40252 19604 40328 19804
use cut_M1M4_1x2 xcut78
transform 1 0 40252 0 1 20564
box 40252 20564 40328 20764
use cut_M1M4_1x2 xcut79
transform 1 0 40252 0 1 21524
box 40252 21524 40328 21724
use cut_M1M4_1x2 xcut80
transform 1 0 40252 0 1 22484
box 40252 22484 40328 22684
use cut_M1M4_1x2 xcut81
transform 1 0 40252 0 1 23444
box 40252 23444 40328 23644
use cut_M1M4_1x2 xcut82
transform 1 0 40252 0 1 24404
box 40252 24404 40328 24604
use cut_M1M4_1x2 xcut83
transform 1 0 40252 0 1 25364
box 40252 25364 40328 25564
use cut_M1M4_1x2 xcut84
transform 1 0 40252 0 1 26324
box 40252 26324 40328 26524
use cut_M1M4_1x2 xcut85
transform 1 0 40252 0 1 27284
box 40252 27284 40328 27484
use cut_M1M4_1x2 xcut86
transform 1 0 40252 0 1 28244
box 40252 28244 40328 28444
use cut_M1M4_1x2 xcut87
transform 1 0 40252 0 1 29204
box 40252 29204 40328 29404
use cut_M1M4_1x2 xcut88
transform 1 0 40252 0 1 30164
box 40252 30164 40328 30364
use cut_M1M4_1x2 xcut89
transform 1 0 40252 0 1 31124
box 40252 31124 40328 31324
use cut_M1M4_1x2 xcut90
transform 1 0 40252 0 1 32084
box 40252 32084 40328 32284
use cut_M1M4_1x2 xcut91
transform 1 0 40252 0 1 33044
box 40252 33044 40328 33244
use cut_M1M4_1x2 xcut92
transform 1 0 40252 0 1 34004
box 40252 34004 40328 34204
use cut_M1M4_1x2 xcut93
transform 1 0 40252 0 1 34964
box 40252 34964 40328 35164
use cut_M1M4_1x2 xcut94
transform 1 0 40252 0 1 35924
box 40252 35924 40328 36124
use cut_M1M4_1x2 xcut95
transform 1 0 40252 0 1 36884
box 40252 36884 40328 37084
use cut_M1M4_1x2 xcut96
transform 1 0 40252 0 1 37844
box 40252 37844 40328 38044
use cut_M1M4_1x2 xcut97
transform 1 0 40252 0 1 38804
box 40252 38804 40328 39004
use cut_M1M4_1x2 xcut98
transform 1 0 40252 0 1 39764
box 40252 39764 40328 39964
use cut_M1M4_1x2 xcut99
transform 1 0 40252 0 1 40724
box 40252 40724 40328 40924
use cut_M1M4_1x2 xcut100
transform 1 0 40252 0 1 41684
box 40252 41684 40328 41884
use cut_M1M4_1x2 xcut101
transform 1 0 40252 0 1 42644
box 40252 42644 40328 42844
use cut_M1M4_1x2 xcut102
transform 1 0 40252 0 1 43604
box 40252 43604 40328 43804
use cut_M1M4_1x2 xcut103
transform 1 0 40252 0 1 44564
box 40252 44564 40328 44764
use cut_M1M4_1x2 xcut104
transform 1 0 40252 0 1 45524
box 40252 45524 40328 45724
use cut_M1M4_1x2 xcut105
transform 1 0 40252 0 1 46484
box 40252 46484 40328 46684
use cut_M1M4_1x2 xcut106
transform 1 0 40252 0 1 47444
box 40252 47444 40328 47644
use cut_M1M4_1x2 xcut107
transform 1 0 40252 0 1 48404
box 40252 48404 40328 48604
<< labels >>
flabel locali s 40252 0 40552 49848 0 FreeSans 400 0 0 0 AVSS
port 2 nsew signal bidirectional
flabel locali s 4516 8558 5092 8778 0 FreeSans 400 0 0 0 VLPFZ
port 1 nsew signal bidirectional
flabel locali s 1060 3882 1636 4102 0 FreeSans 400 0 0 0 VLPF
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 40552 49848
<< end >>
