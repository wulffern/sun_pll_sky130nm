magic
tech sky130B
magscale 1 2
timestamp 1679853665
<< locali >>
rect 0 5696 4344 5936
rect 0 240 240 5696
rect 384 5312 3960 5552
rect 384 624 624 5312
rect 1200 4786 1428 4846
rect 1632 4698 2064 4758
rect 1632 4346 1860 4406
rect 1800 4230 1860 4346
rect 1632 4170 1860 4230
rect 1170 914 1230 2734
rect 2004 2646 2064 4698
rect 1632 2586 2064 2646
rect 2004 886 2064 2586
rect 3180 2234 3612 2294
rect 3180 1882 3408 1942
rect 3348 1766 3408 1882
rect 3180 1706 3408 1766
rect 3552 1414 3612 2234
rect 3180 1354 3612 1414
rect 3552 886 3612 1354
rect 1632 826 2064 886
rect 3180 826 3612 886
rect 3720 624 3960 5312
rect 384 384 3960 624
rect 4104 240 4344 5696
rect 0 0 4344 240
<< metal1 >>
rect 1632 4874 1860 4934
rect 1632 4522 3408 4582
rect 3348 2470 3408 4522
rect 1632 2410 2976 2470
rect 3180 2410 3408 2470
rect 2916 1502 2976 2410
rect 3348 2118 3408 2410
rect 3180 2058 3408 2118
rect 2748 1442 2976 1502
rect 2916 1238 2976 1442
rect 2916 1178 3180 1238
rect 660 384 876 988
rect 1524 384 1740 886
rect 2208 0 2424 988
rect 2916 974 2976 1178
rect 2748 914 2976 974
rect 3072 0 3288 886
<< metal2 >>
rect 1632 4934 4236 4950
rect 1632 4874 4344 4934
rect 108 4846 1200 4862
rect 0 4786 1200 4846
rect 1632 4582 4236 4598
rect 1632 4522 4344 4582
rect 108 4494 1200 4510
rect 0 4434 1200 4494
rect 108 2382 2576 2398
rect 0 2368 2576 2382
rect 0 2322 2748 2368
rect 2500 2292 2748 2322
rect 108 2030 2748 2046
rect 0 1970 2748 2030
rect 108 974 1200 990
rect 0 914 1200 974
use cut_M1M2_2x1  cut_M1M2_2x1_0
timestamp 1677625200
transform 1 0 1524 0 1 4874
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_1
timestamp 1677625200
transform 1 0 3072 0 1 2410
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_2
timestamp 1677625200
transform 1 0 1524 0 1 4522
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_3
timestamp 1677625200
transform 1 0 3072 0 1 2058
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_4
timestamp 1677625200
transform 1 0 2640 0 1 1442
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_5
timestamp 1677625200
transform 1 0 1524 0 1 2410
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_6
timestamp 1677625200
transform 1 0 3072 0 1 1178
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_7
timestamp 1677625200
transform 1 0 2640 0 1 914
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_8
timestamp 1677625200
transform 1 0 2224 0 1 0
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_9
timestamp 1677625200
transform 1 0 2224 0 1 900
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_10
timestamp 1677625200
transform 1 0 3088 0 1 0
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_11
timestamp 1677625200
transform 1 0 3088 0 1 826
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_12
timestamp 1677625200
transform 1 0 676 0 1 384
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_13
timestamp 1677625200
transform 1 0 676 0 1 900
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_14
timestamp 1677625200
transform 1 0 1540 0 1 384
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_15
timestamp 1677625200
transform 1 0 1540 0 1 826
box 0 0 184 68
use cut_M1M3_2x1  cut_M1M3_2x1_0
timestamp 1677625200
transform 1 0 1108 0 1 4434
box 0 0 200 76
use cut_M1M3_2x1  cut_M1M3_2x1_1
timestamp 1677625200
transform 1 0 2656 0 1 1970
box 0 0 200 76
use cut_M1M3_2x1  cut_M1M3_2x1_2
timestamp 1677625200
transform 1 0 1524 0 1 4874
box 0 0 200 76
use cut_M1M3_2x1  cut_M1M3_2x1_3
timestamp 1677625200
transform 1 0 1524 0 1 4522
box 0 0 200 76
use cut_M1M3_2x1  cut_M1M3_2x1_4
timestamp 1677625200
transform 1 0 1108 0 1 914
box 0 0 200 76
use cut_M1M3_2x1  cut_M1M3_2x1_5
timestamp 1677625200
transform 1 0 1108 0 1 4786
box 0 0 200 76
use cut_M1M3_2x1  cut_M1M3_2x1_6
timestamp 1677625200
transform 1 0 2656 0 1 2284
box 0 0 200 76
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM#0  xa1 ../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1679853665
transform 1 0 768 0 1 768
box -180 -132 1260 1892
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM#0  xa2
timestamp 1679853665
transform 1 0 768 0 1 2528
box -180 -132 1260 1892
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL#0  xa3 ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 0
transform 1 0 768 0 1 4288
box 0 0 1 1
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLA#0  xa4 ../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1679853665
transform 1 0 768 0 1 4640
box -180 -132 1260 660
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLCM  xb1 ../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1679853665
transform -1 0 3576 0 1 768
box 0 -132 1440 660
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDLCM  xb2
timestamp 1679853665
transform -1 0 3576 0 1 1296
box 0 -132 1440 660
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL#0  xb3 ../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1677625200
transform -1 0 3576 0 1 1824
box 0 -132 1440 484
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_PCHDL#0  xb4
timestamp 1677625200
transform -1 0 3576 0 1 2176
box 0 -132 1440 484
<< labels >>
flabel locali s 3720 384 3960 5552 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
flabel locali s 4104 0 4344 5936 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel metal2 s 0 1970 216 2030 0 FreeSans 400 0 0 0 CP_UP_N
port 2 nsew
flabel metal2 s 4128 4522 4344 4582 0 FreeSans 400 0 0 0 LPF
port 3 nsew
flabel metal2 s 0 4434 216 4494 0 FreeSans 400 0 0 0 CP_DOWN
port 4 nsew
flabel metal2 s 0 914 216 974 0 FreeSans 400 0 0 0 VBN
port 5 nsew
flabel metal2 s 4128 4874 4344 4934 0 FreeSans 400 0 0 0 LPFZ
port 7 nsew
flabel metal2 s 0 2322 216 2382 0 FreeSans 400 0 0 0 PWRUP_1V8
port 8 nsew
flabel metal2 s 0 4786 216 4846 0 FreeSans 400 0 0 0 KICK
port 9 nsew
<< end >>
