magic
tech sky130B
magscale 1 1
timestamp 1720908000
<< checkpaint >>
rect 0 0 1014 1440
<< locali >>
rect 894 0 1014 1440
rect 0 0 1014 120
rect 0 1320 1014 1440
rect 0 0 120 1440
rect 894 0 1014 1440
rect 408 265 492 295
rect 492 265 522 295
rect 510 339 600 369
rect 510 1189 624 1219
rect 408 441 510 471
rect 510 339 540 1219
rect 570 309 624 339
rect 678 221 1014 251
rect 678 397 1014 427
rect 0 258 138 288
rect 0 434 138 464
<< m2 >>
rect 906 309 1014 339
rect 0 265 108 295
rect 906 309 1014 339
rect 500 309 624 347
rect 500 309 960 347
rect 500 309 538 347
rect 0 265 108 295
rect 284 265 408 303
rect 54 265 284 303
rect 284 265 322 303
use SUNTR_NCHDL xa2 ../SUN_TR_SKY130NM
transform 1 0 192 0 1 192
box 192 192 822 368
use SUNTR_NCHDLCM xa3 ../SUN_TR_SKY130NM
transform 1 0 192 0 1 368
box 192 368 822 1248
use cut_M1M3_2x1 xcut0 
transform 1 0 578 0 1 309
box 578 309 678 347
use cut_M1M3_2x1 xcut1 
transform 1 0 362 0 1 265
box 362 265 462 303
<< labels >>
flabel locali s 894 0 1014 1440 0 FreeSans 400 0 0 0 AVSS
port 3 nsew signal bidirectional
flabel m2 s 906 309 1014 339 0 FreeSans 400 0 0 0 IBPSR_1U
port 1 nsew signal bidirectional
flabel m2 s 0 265 108 295 0 FreeSans 400 0 0 0 PWRUP_1V8_N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1014 1440
<< end >>
