magic
tech sky130B
magscale 1 2
timestamp 1679853665
<< locali >>
rect 0 2640 2028 2880
rect 0 928 240 2640
rect 1020 2378 1248 2438
rect 1020 942 1080 2378
rect 0 868 276 928
rect 816 882 1080 942
rect 0 576 240 868
rect 1020 738 1080 882
rect 1788 854 2028 2640
rect 1356 794 2028 854
rect 1020 678 1200 738
rect 1140 618 1248 678
rect 0 516 276 576
rect 816 530 1044 590
rect 0 240 240 516
rect 1788 502 2028 794
rect 1356 442 2028 502
rect 1788 240 2028 442
rect 0 0 2028 240
<< metal2 >>
rect 1000 678 1920 694
rect 1000 618 2028 678
rect 108 590 816 606
rect 0 530 816 590
use cut_M1M3_2x1  cut_M1M3_2x1_0
timestamp 1677625200
transform 1 0 724 0 1 530
box 0 0 200 76
use cut_M1M3_2x1  cut_M1M3_2x1_1
timestamp 1677625200
transform 1 0 1156 0 1 618
box 0 0 200 76
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDL#1  xa2 ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 0
transform 1 0 384 0 1 384
box 0 0 1 1
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NCHDLCM#1  xa3 ../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1677625200
transform 1 0 384 0 1 736
box -180 -132 1260 1892
<< labels >>
flabel locali s 1788 0 2028 2880 0 FreeSans 400 0 0 0 AVSS
port 3 nsew
flabel metal2 s 1812 618 2028 678 0 FreeSans 400 0 0 0 IBPSR_1U
port 1 nsew
flabel metal2 s 0 530 216 590 0 FreeSans 400 0 0 0 PWRUP_1V8_N
port 2 nsew
<< end >>
