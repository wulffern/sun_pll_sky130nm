magic
tech sky130B
magscale 1 2
timestamp 1681509600
<< checkpaint >>
rect 0 0 33680 960
<< m1 >>
rect 120 -40 33640 40
rect 33560 40 33640 120
rect 120 120 33480 200
rect 33560 120 33640 200
rect 120 200 200 280
rect 33560 200 33640 280
rect 120 280 200 360
rect 280 280 33640 360
rect 120 360 200 440
rect 33560 360 33640 440
rect 120 440 33480 520
rect 33560 440 33640 520
rect 120 520 200 600
rect 33560 520 33640 600
rect 120 600 200 680
rect 280 600 33640 680
rect 120 680 200 760
rect 120 760 33640 840
<< m2 >>
rect 120 -40 33640 40
rect 33560 40 33640 120
rect 120 120 33480 200
rect 33560 120 33640 200
rect 120 200 200 280
rect 33560 200 33640 280
rect 120 280 200 360
rect 280 280 33640 360
rect 120 360 200 440
rect 33560 360 33640 440
rect 120 440 33480 520
rect 33560 440 33640 520
rect 120 520 200 600
rect 33560 520 33640 600
rect 120 600 200 680
rect 280 600 33640 680
rect 120 680 200 760
rect 120 760 33640 840
<< locali >>
rect 120 -40 33640 40
rect 33560 40 33640 120
rect 120 120 33480 200
rect 33560 120 33640 200
rect 120 200 200 280
rect 33560 200 33640 280
rect 120 280 200 360
rect 280 280 33640 360
rect 120 360 200 440
rect 33560 360 33640 440
rect 120 440 33480 520
rect 33560 440 33640 520
rect 120 520 200 600
rect 33560 520 33640 600
rect 120 600 200 680
rect 280 600 33640 680
rect 120 680 200 760
rect 120 760 33640 840
<< v1 >>
rect 33160 -28 33400 28
rect 280 132 520 188
rect 33160 292 33400 348
rect 280 452 520 508
rect 33160 612 33400 668
rect 280 772 520 828
<< v2 >>
rect 33160 -32 33400 32
rect 280 128 520 192
rect 33160 288 33400 352
rect 280 448 520 512
rect 33160 608 33400 672
rect 280 768 520 832
<< viali >>
rect 33160 -28 33400 28
rect 280 132 520 188
rect 33160 292 33400 348
rect 280 452 520 508
rect 33160 612 33400 668
rect 280 772 520 828
<< m3 >>
rect 120 -40 33640 40
rect 120 -40 33640 40
rect 33560 40 33640 120
rect 120 120 33240 200
rect 33320 120 33480 200
rect 33560 120 33640 200
rect 120 200 200 280
rect 33560 200 33640 280
rect 120 280 200 360
rect 280 280 360 360
rect 440 280 33640 360
rect 120 360 200 440
rect 33560 360 33640 440
rect 120 440 33480 520
rect 33560 440 33640 520
rect 120 520 200 600
rect 33560 520 33640 600
rect 120 600 200 680
rect 280 600 33640 680
rect 120 680 200 760
rect 120 760 33640 840
rect 120 760 33640 840
<< rm3 >>
rect 33240 120 33320 200
rect 360 280 440 360
<< labels >>
flabel m3 s 120 -40 33640 40 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel m3 s 120 760 33640 840 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 33680 960
<< end >>
