magic
tech sky130B
magscale 1 1
timestamp 1720908000
<< checkpaint >>
rect 0 0 16840 480
<< m1 >>
rect 60 -20 16820 20
rect 16780 20 16820 60
rect 60 60 16740 100
rect 16780 60 16820 100
rect 60 100 100 140
rect 16780 100 16820 140
rect 60 140 100 180
rect 140 140 16820 180
rect 60 180 100 220
rect 16780 180 16820 220
rect 60 220 16740 260
rect 16780 220 16820 260
rect 60 260 100 300
rect 16780 260 16820 300
rect 60 300 100 340
rect 140 300 16820 340
rect 60 340 100 380
rect 60 380 16820 420
<< m2 >>
rect 60 -20 16820 20
rect 16780 20 16820 60
rect 60 60 16740 100
rect 16780 60 16820 100
rect 60 100 100 140
rect 16780 100 16820 140
rect 60 140 100 180
rect 140 140 16820 180
rect 60 180 100 220
rect 16780 180 16820 220
rect 60 220 16740 260
rect 16780 220 16820 260
rect 60 260 100 300
rect 16780 260 16820 300
rect 60 300 100 340
rect 140 300 16820 340
rect 60 340 100 380
rect 60 380 16820 420
<< locali >>
rect 60 -20 16820 20
rect 16780 20 16820 60
rect 60 60 16740 100
rect 16780 60 16820 100
rect 60 100 100 140
rect 16780 100 16820 140
rect 60 140 100 180
rect 140 140 16820 180
rect 60 180 100 220
rect 16780 180 16820 220
rect 60 220 16740 260
rect 16780 220 16820 260
rect 60 260 100 300
rect 16780 260 16820 300
rect 60 300 100 340
rect 140 300 16820 340
rect 60 340 100 380
rect 60 380 16820 420
<< v1 >>
rect 16580 -14 16700 14
rect 140 66 260 94
rect 16580 146 16700 174
rect 140 226 260 254
rect 16580 306 16700 334
rect 140 386 260 414
<< v2 >>
rect 16580 -16 16700 16
rect 140 64 260 96
rect 16580 144 16700 176
rect 140 224 260 256
rect 16580 304 16700 336
rect 140 384 260 416
<< viali >>
rect 16580 -14 16700 14
rect 140 66 260 94
rect 16580 146 16700 174
rect 140 226 260 254
rect 16580 306 16700 334
rect 140 386 260 414
<< m3 >>
rect 60 -20 16820 20
rect 60 -20 16820 20
rect 16780 20 16820 60
rect 60 60 16620 100
rect 16660 60 16740 100
rect 16780 60 16820 100
rect 60 100 100 140
rect 16780 100 16820 140
rect 60 140 100 180
rect 140 140 180 180
rect 220 140 16820 180
rect 60 180 100 220
rect 16780 180 16820 220
rect 60 220 16740 260
rect 16780 220 16820 260
rect 60 260 100 300
rect 16780 260 16820 300
rect 60 300 100 340
rect 140 300 16820 340
rect 60 340 100 380
rect 60 380 16820 420
rect 60 380 16820 420
<< rm3 >>
rect 16620 60 16660 100
rect 180 140 220 180
<< labels >>
flabel m3 s 60 -20 16820 20 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel m3 s 60 380 16820 420 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 16840 480
<< end >>
