magic
tech sky130B
magscale 1 2
timestamp 1681511206
<< locali >>
rect 24003 68549 24658 69221
rect 24003 67906 24009 68549
rect 24652 67906 24658 68549
rect 24003 67900 24658 67906
rect -2000 66676 35028 67000
rect -2000 66448 34426 66676
rect 34654 66448 35028 66676
rect -2000 66000 35028 66448
rect 2080 64696 2320 66000
rect -1772 63760 -1760 63880
rect 3600 59368 3840 66000
rect 17060 64972 17300 66000
rect 31008 65168 31248 66000
rect 1816 57480 2056 59120
rect 4818 55655 4878 55726
rect 5680 55014 6120 55020
rect 5680 54786 5686 55014
rect 5914 54786 6120 55014
rect 5680 54780 6120 54786
rect 5388 53780 5680 54020
rect 5388 51000 5628 51520
rect -2000 50976 24003 51000
rect 24658 50976 39000 51000
rect -2000 50569 39000 50976
rect -2000 50414 14706 50569
rect -2000 50186 1386 50414
rect 1614 50336 14706 50414
rect 14939 50336 39000 50569
rect 1614 50268 39000 50336
rect 1614 50186 29850 50268
rect -2000 50064 29850 50186
rect 30054 50064 39000 50268
rect -2000 50000 39000 50064
<< viali >>
rect 24009 67906 24652 68549
rect 34426 66448 34654 66676
rect 29060 60392 29288 60620
rect 5566 59106 5611 59151
rect 25010 58962 25074 59026
rect 34420 58576 34660 58816
rect 29054 58192 29294 58432
rect 5656 55754 5716 55814
rect 4818 55595 4878 55655
rect 5686 54786 5914 55014
rect 5680 53780 5920 54020
rect 1380 52384 1620 52624
rect 14714 52424 14900 52578
rect 24003 50976 24658 51631
rect 1386 50186 1614 50414
rect 14706 50336 14939 50569
rect 29850 50064 30054 50268
<< metal1 >>
rect -1128 78014 -1056 78020
rect -1321 73395 -1250 73428
rect -1327 73324 -1321 73395
rect -1250 73324 -1244 73395
rect -1321 67328 -1250 73324
rect -1128 67542 -1056 77942
rect 2554 78014 2626 78020
rect 2554 77596 2626 77942
rect 24003 68549 24658 68561
rect 24003 67906 24009 68549
rect 24652 67906 24658 68549
rect -1128 67464 -1056 67470
rect 2896 67542 2968 67548
rect 2640 67328 2711 67334
rect -1327 67257 -1321 67328
rect -1250 67257 -1244 67328
rect -1986 65300 -1980 65420
rect -1860 65300 -1854 65420
rect -1980 63892 -1860 65300
rect -1980 63766 -1860 63772
rect 2640 63590 2711 67257
rect 2896 63944 2968 67470
rect 8184 67328 8255 67334
rect 5511 65420 5654 65445
rect 5511 65300 5520 65420
rect 5640 65300 5654 65420
rect 5511 65243 5654 65300
rect 2896 63866 2968 63872
rect 2640 63513 2711 63519
rect -1708 61398 -1602 61417
rect -1708 61322 -1695 61398
rect -1619 61322 -1602 61398
rect -1708 61307 -1602 61322
rect -1996 59914 -1990 59974
rect -1930 59914 -1924 59974
rect -1990 58810 -1930 59914
rect -1990 58744 -1930 58750
rect -1695 56663 -1619 61307
rect 5560 59151 5617 65243
rect 5560 59106 5566 59151
rect 5611 59106 5617 59151
rect 5560 59094 5617 59106
rect 3411 58809 3471 58815
rect -1695 56587 -1444 56663
rect -1672 56146 -1612 56152
rect -1672 51224 -1612 56086
rect -1520 51575 -1444 56587
rect 3161 55814 3221 55820
rect 2866 55655 2926 55661
rect 1368 52624 1632 52630
rect 1368 52384 1380 52624
rect 1620 52384 1632 52624
rect 1368 52378 1632 52384
rect -1520 51493 -1444 51499
rect -1678 51164 -1672 51224
rect -1612 51164 -1606 51224
rect 1380 50414 1620 52378
rect 2293 51990 2299 52050
rect 2359 51990 2365 52050
rect 2299 51769 2359 51990
rect 2299 51703 2359 51709
rect 2866 51559 2926 55595
rect 3161 51788 3221 55754
rect 3411 54268 3471 58749
rect 5626 55820 5748 55858
rect 5626 55748 5650 55820
rect 5722 55748 5748 55820
rect 5626 55695 5748 55748
rect 4806 55589 4812 55661
rect 4872 55655 4890 55661
rect 4878 55595 4890 55655
rect 4872 55589 4890 55595
rect 8184 55270 8255 67257
rect 8184 55193 8255 55199
rect 23818 59212 23878 59218
rect 5680 55014 5920 55026
rect 5680 54786 5686 55014
rect 5914 54786 5920 55014
rect 3411 54202 3471 54208
rect 5445 54268 5505 54274
rect 5445 51878 5505 54208
rect 5680 54032 5920 54786
rect 5674 54020 5926 54032
rect 5674 53780 5680 54020
rect 5920 53780 5926 54020
rect 5674 53768 5926 53780
rect 7313 52967 7372 52973
rect 7313 51884 7372 52908
rect 14678 52578 14944 52624
rect 14678 52424 14714 52578
rect 14900 52489 14944 52578
rect 14900 52424 14945 52489
rect 14678 52384 14945 52424
rect 14680 52308 14945 52384
rect 7756 51984 7762 52060
rect 7838 51984 7844 52060
rect 5445 51812 5505 51818
rect 7312 51878 7372 51884
rect 7312 51812 7372 51818
rect 3161 51722 3221 51728
rect 7762 51572 7838 51984
rect 8118 51624 8178 51630
rect 2866 51493 2926 51499
rect 7756 51496 7762 51572
rect 7838 51496 7844 51572
rect 8118 51224 8178 51564
rect 8118 51158 8178 51164
rect 1380 50186 1386 50414
rect 1614 50186 1620 50414
rect 14700 50569 14945 52308
rect 23818 51624 23878 59152
rect 24003 51637 24658 67906
rect 34420 66676 34660 66688
rect 34420 66448 34426 66676
rect 34654 66448 34660 66676
rect 32022 65408 32082 65414
rect 26762 65348 27060 65408
rect 27120 65348 27126 65408
rect 29054 60620 29294 60632
rect 29054 60392 29060 60620
rect 29288 60392 29294 60620
rect 26404 59212 26464 59218
rect 25004 59026 25080 59038
rect 25004 58962 25010 59026
rect 25074 58962 25080 59026
rect 25004 52060 25080 58962
rect 26404 58828 26464 59152
rect 29054 58438 29294 60392
rect 30346 58970 30406 60060
rect 32022 59486 32082 65348
rect 32022 59420 32082 59426
rect 34420 58838 34660 66448
rect 38670 59426 38676 59486
rect 38736 59426 38742 59486
rect 34388 58816 34702 58838
rect 34388 58576 34420 58816
rect 34660 58576 34702 58816
rect 34388 58552 34702 58576
rect 29042 58432 29306 58438
rect 29042 58192 29054 58432
rect 29294 58192 29306 58432
rect 29042 58186 29306 58192
rect 24998 51984 25004 52060
rect 25080 51984 25086 52060
rect 36260 51922 36320 52054
rect 38676 51922 38736 59426
rect 38670 51862 38676 51922
rect 38736 51862 38742 51922
rect 36260 51856 36320 51862
rect 23818 51558 23878 51564
rect 23991 51631 24670 51637
rect 23991 50976 24003 51631
rect 24658 50976 24670 51631
rect 23991 50970 24670 50976
rect 14700 50336 14706 50569
rect 14939 50336 14945 50569
rect 14700 50324 14945 50336
rect 29844 50274 30060 50280
rect 1380 50174 1620 50186
rect 29838 50058 29844 50274
rect 30060 50058 30066 50274
rect 29844 50052 30060 50058
<< via1 >>
rect -1128 77942 -1056 78014
rect -1321 73324 -1250 73395
rect 2554 77942 2626 78014
rect -1128 67470 -1056 67542
rect 2896 67470 2968 67542
rect -1321 67257 -1250 67328
rect 2640 67257 2711 67328
rect -1980 65300 -1860 65420
rect -1980 63772 -1860 63892
rect 8184 67257 8255 67328
rect 5520 65300 5640 65420
rect 2896 63872 2968 63944
rect 2640 63519 2711 63590
rect -1695 61322 -1619 61398
rect -1990 59914 -1930 59974
rect -1990 58750 -1930 58810
rect 3411 58749 3471 58809
rect -1672 56086 -1612 56146
rect 3161 55754 3221 55814
rect 2866 55595 2926 55655
rect -1520 51499 -1444 51575
rect -1672 51164 -1612 51224
rect 2299 51990 2359 52050
rect 2299 51709 2359 51769
rect 5650 55814 5722 55820
rect 5650 55754 5656 55814
rect 5656 55754 5716 55814
rect 5716 55754 5722 55814
rect 5650 55748 5722 55754
rect 4812 55655 4872 55661
rect 4812 55595 4818 55655
rect 4818 55595 4872 55655
rect 4812 55589 4872 55595
rect 8184 55199 8255 55270
rect 23818 59152 23878 59212
rect 3411 54208 3471 54268
rect 5445 54208 5505 54268
rect 7313 52908 7372 52967
rect 7762 51984 7838 52060
rect 5445 51818 5505 51878
rect 7312 51818 7372 51878
rect 3161 51728 3221 51788
rect 2866 51499 2926 51559
rect 7762 51496 7838 51572
rect 8118 51564 8178 51624
rect 8118 51164 8178 51224
rect 27060 65348 27120 65408
rect 32022 65348 32082 65408
rect 26404 59152 26464 59212
rect 32022 59426 32082 59486
rect 38676 59426 38736 59486
rect 25004 51984 25080 52060
rect 36260 51862 36320 51922
rect 38676 51862 38736 51922
rect 23818 51564 23878 51624
rect 29844 50268 30060 50274
rect 29844 50064 29850 50268
rect 29850 50064 30054 50268
rect 30054 50064 30060 50268
rect 29844 50058 30060 50064
<< metal2 >>
rect -1134 77942 -1128 78014
rect -1056 77942 2554 78014
rect 2626 77942 2632 78014
rect -1321 73395 -1250 73401
rect -1250 73324 2645 73395
rect -1321 73318 -1250 73324
rect 2574 72919 2645 73324
rect -1134 67470 -1128 67542
rect -1056 67470 2896 67542
rect 2968 67470 2974 67542
rect -1321 67328 -1250 67334
rect -1250 67257 2640 67328
rect 2711 67257 8184 67328
rect 8255 67257 8261 67328
rect -1321 67251 -1250 67257
rect 11938 65739 29268 65744
rect 11938 65533 29057 65739
rect 29263 65533 29272 65739
rect 11938 65528 29268 65533
rect -1980 65420 -1860 65426
rect -1860 65300 5520 65420
rect 5640 65300 5646 65420
rect 12098 65340 12314 65528
rect 27060 65408 27120 65414
rect 27120 65348 32022 65408
rect 32082 65348 32088 65408
rect 27060 65342 27120 65348
rect -1980 65294 -1860 65300
rect 10029 65124 10038 65340
rect 10254 65124 12314 65340
rect -1986 63772 -1980 63892
rect -1860 63772 -1854 63892
rect 2096 63872 2896 63944
rect 2968 63872 2974 63944
rect 2099 63519 2640 63590
rect 2711 63519 2717 63590
rect -1957 63432 -1948 63488
rect -1892 63432 -1883 63488
rect -1708 61398 -1602 61417
rect -1708 61322 -1695 61398
rect -1619 61322 -1602 61398
rect -1708 61307 -1602 61322
rect -2100 61028 -1730 61030
rect -2107 60972 -2098 61028
rect -2042 60972 -1730 61028
rect -2100 60970 -1730 60972
rect -1990 59974 -1930 59980
rect -1990 59908 -1930 59914
rect 38676 59486 38736 59492
rect 32016 59426 32022 59486
rect 32082 59426 38676 59486
rect 38736 59426 39156 59486
rect 38676 59420 38736 59426
rect 23812 59152 23818 59212
rect 23878 59152 26404 59212
rect 26464 59152 26470 59212
rect -1996 58750 -1990 58810
rect -1930 58809 3790 58810
rect -1930 58750 3411 58809
rect 3405 58749 3411 58750
rect 3471 58750 3790 58809
rect 3471 58749 3477 58750
rect 2392 58230 2448 58237
rect -2109 58170 -2100 58230
rect -2040 58228 2450 58230
rect -2040 58172 2392 58228
rect 2448 58172 2450 58228
rect -2040 58170 2450 58172
rect 2392 58163 2448 58170
rect -1959 58030 -1950 58090
rect -1890 58088 2230 58090
rect -1890 58032 2172 58088
rect 2228 58032 2237 58088
rect -1890 58030 2230 58032
rect 1996 56874 2170 56934
rect 2230 56874 2239 56934
rect -1678 56086 -1672 56146
rect -1612 56086 -1606 56146
rect 5626 55820 5748 55858
rect 5626 55814 5650 55820
rect 3155 55754 3161 55814
rect 3221 55754 5650 55814
rect 5626 55748 5650 55754
rect 5722 55748 5748 55820
rect 5626 55695 5748 55748
rect 4812 55661 4872 55667
rect 2860 55595 2866 55655
rect 2926 55595 4812 55655
rect 4812 55583 4872 55589
rect 8178 55199 8184 55270
rect 8255 55199 9243 55270
rect 1996 54762 2390 54822
rect 2450 54762 2459 54822
rect 3405 54208 3411 54268
rect 3471 54208 5445 54268
rect 5505 54208 5511 54268
rect -2132 53618 -1560 53694
rect 7307 52908 7313 52967
rect 7372 52908 9077 52967
rect 7762 52060 7838 52066
rect 25004 52060 25080 52066
rect 2299 52050 2359 52056
rect 2359 51990 5926 52050
rect 2299 51984 2359 51990
rect 5866 51878 5926 51990
rect 7838 51984 11172 52060
rect 7762 51978 7838 51984
rect 11096 51892 11172 51984
rect 12502 51984 25004 52060
rect 12502 51892 12578 51984
rect 25004 51978 25080 51984
rect 38676 51922 38736 51928
rect 5439 51818 5445 51878
rect 5505 51818 7312 51878
rect 7372 51818 7378 51878
rect 11096 51816 12578 51892
rect 36254 51862 36260 51922
rect 36320 51862 38676 51922
rect 38676 51856 38736 51862
rect -2136 51709 2299 51769
rect 2359 51709 2365 51769
rect 3155 51728 3161 51788
rect 3221 51728 4127 51788
rect -1526 51572 -1520 51575
rect -2133 51499 -1520 51572
rect -1444 51572 -1438 51575
rect 7762 51572 7838 51578
rect -1444 51559 7762 51572
rect -1444 51499 2866 51559
rect 2926 51499 7762 51559
rect -2133 51496 7762 51499
rect 8112 51564 8118 51624
rect 8178 51564 23818 51624
rect 23878 51564 23884 51624
rect 7762 51490 7838 51496
rect -1672 51224 -1612 51230
rect -1612 51164 8118 51224
rect 8178 51164 8184 51224
rect -1672 51158 -1612 51164
rect 29844 50274 30060 50280
rect 29840 50063 29844 50269
rect 30060 50063 30064 50269
rect 29844 50052 30060 50058
<< via2 >>
rect 29057 65533 29263 65739
rect 10038 65124 10254 65340
rect -1948 63432 -1892 63488
rect -2098 60972 -2042 61028
rect -2100 58170 -2040 58230
rect 2392 58172 2448 58228
rect -1950 58030 -1890 58090
rect 2172 58032 2228 58088
rect 2170 56874 2230 56934
rect 2390 54762 2450 54822
rect 29849 50063 30055 50269
<< metal3 >>
rect 29052 65739 29268 65744
rect 29052 65533 29057 65739
rect 29263 65533 29268 65739
rect 10033 65340 10259 65345
rect 10033 65124 10038 65340
rect 10254 65124 10259 65340
rect 29052 65192 29268 65533
rect 10033 65119 10259 65124
rect -1953 63488 -1887 63493
rect -1953 63432 -1948 63488
rect -1892 63432 -1887 63488
rect -1953 63427 -1887 63432
rect -2103 61028 -2037 61033
rect -2103 60972 -2098 61028
rect -2042 60972 -2037 61028
rect -2103 60967 -2037 60972
rect -2100 58235 -2040 60967
rect -2105 58230 -2035 58235
rect -2105 58170 -2100 58230
rect -2040 58170 -2035 58230
rect -2105 58165 -2035 58170
rect -1950 58095 -1890 63427
rect 2387 58228 2453 58233
rect 2387 58172 2392 58228
rect 2448 58172 2453 58228
rect 2387 58167 2453 58172
rect -1955 58090 -1885 58095
rect -1955 58030 -1950 58090
rect -1890 58030 -1885 58090
rect -1955 58025 -1885 58030
rect 2167 58088 2233 58093
rect 2167 58032 2172 58088
rect 2228 58032 2233 58088
rect 2167 58027 2233 58032
rect 2170 56939 2230 58027
rect 2165 56934 2235 56939
rect 2165 56874 2170 56934
rect 2230 56874 2235 56934
rect 2165 56869 2235 56874
rect 2390 54827 2450 58167
rect 2385 54822 2455 54827
rect 2385 54762 2390 54822
rect 2450 54762 2455 54822
rect 2385 54757 2455 54762
rect 29844 50269 30060 52796
rect 29844 50063 29849 50269
rect 30055 50063 30060 50269
rect 29844 50058 30060 50063
use SUN_PLL_PFD  xaa0
timestamp 1681511206
transform 1 0 -2000 0 1 52000
box 0 0 4056 5760
use SUN_PLL_CP  xaa1
timestamp 1681511206
transform 1 0 -2000 0 1 59000
box 0 0 4344 5936
use SUN_PLL_KICK  xaa3
timestamp 1681511206
transform 1 0 3600 0 1 54400
box 0 0 4128 5936
use SUN_PLL_BUF  xaa4
timestamp 1681511206
transform 1 0 9000 0 1 52000
box 0 0 14784 13184
use SUN_PLL_ROSC  xaa5
timestamp 1681511206
transform 1 0 25000 0 1 60000
box 0 0 6576 5408
use SUN_PLL_DIVN  xaa6
timestamp 1681511206
transform 1 0 25000 0 1 52000
box 0 0 14136 7036
use SUN_PLL_LPF  xbb0
timestamp 1681511206
transform 1 0 -2000 0 1 69000
box 0 0 40552 24888
use SUN_PLL_BIAS  xbb1
timestamp 1681511206
transform 1 0 3600 0 1 51200
box 0 0 2028 2880
<< labels >>
flabel locali -1962 66042 -732 66844 0 FreeSans 1600 0 0 0 AVDD
port 0 nsew
flabel locali -1808 50056 -578 50858 0 FreeSans 1600 0 0 0 AVSS
port 1 nsew
flabel metal2 -2133 51496 -2057 51572 0 FreeSans 800 0 0 0 PWRUP_1V8
port 2 nsew
flabel metal2 -2132 53618 -2056 53694 0 FreeSans 800 0 0 0 CK_REF
port 3 nsew
flabel metal2 39096 59426 39156 59486 0 FreeSans 800 0 0 0 CK
port 4 nsew
flabel metal2 -2136 51709 -2076 51769 0 FreeSans 800 0 0 0 IBPSR_1U
port 5 nsew
flabel metal1 -1128 67542 -1056 73256 0 FreeSans 800 0 0 0 VLPZ
flabel space 9670 65528 29057 65744 0 FreeSans 800 0 0 0 VDD_ROSC
flabel metal2 -1250 67257 2640 67328 0 FreeSans 800 0 0 0 VLPF
<< end >>
