magic
tech sky130B
magscale 1 2
timestamp 1667257200
<< checkpaint >>
rect 0 0 39832 22068
<< locali >>
rect 39532 0 39832 22068
rect 0 0 39832 300
rect 0 21768 39832 22068
rect 0 0 300 22068
rect 39532 0 39832 22068
rect 300 460 460 572
rect 300 4696 460 4808
rect 300 8932 460 9044
rect 300 13168 460 13280
rect 300 17404 460 17516
rect 4516 20826 5092 21046
rect 1060 3882 1636 4102
<< m3 >>
rect 22400 0 22616 484
rect 39268 404 39608 480
rect 39268 1364 39608 1440
rect 39268 2324 39608 2400
<< m1 >>
rect 1152 8118 1364 8178
rect 1364 3882 4608 3942
rect 1364 3882 1424 8178
rect 1152 16590 1508 16650
rect 1508 12354 4608 12414
rect 1508 12354 1568 16650
rect 4608 20826 4760 20886
rect 4760 3124 5848 3184
rect 4760 3124 4820 20886
<< m2 >>
rect 1160 12354 1388 12430
rect 1388 8118 4616 8194
rect 1388 8118 1464 12430
rect 1160 20826 1676 20902
rect 1676 16590 4616 16666
rect 1676 16590 1752 20902
rect 1160 3882 1324 3958
rect 1324 1204 5848 1280
rect 1324 2164 5848 2240
rect 1324 1204 1400 3958
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8 xa1
transform 1 0 444 0 1 444
box 444 444 5708 4680
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8 xa2
transform 1 0 444 0 1 4680
box 444 4680 5708 8916
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8 xa3
transform 1 0 444 0 1 8916
box 444 8916 5708 13152
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8 xa4
transform 1 0 444 0 1 13152
box 444 13152 5708 17388
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_RPPO8 xa5
transform 1 0 444 0 1 17388
box 444 17388 5708 21624
use CAP_LPF xb1
transform -1 0 39388 0 1 444
box 39388 444 73068 1404
use CAP_LPF xb2
transform -1 0 39388 0 1 1404
box 39388 1404 73068 2364
use CAP_LPF xb3
transform -1 0 39388 0 1 2364
box 39388 2364 73068 3324
use cut_M1M4_2x1 
transform 1 0 22408 0 1 0
box 22408 0 22608 76
use cut_M1M2_2x1 
transform 1 0 1060 0 1 8118
box 1060 8118 1244 8186
use cut_M1M2_2x1 
transform 1 0 4516 0 1 3882
box 4516 3882 4700 3950
use cut_M1M3_2x1 
transform 1 0 1060 0 1 12354
box 1060 12354 1260 12430
use cut_M1M3_2x1 
transform 1 0 4516 0 1 8118
box 4516 8118 4716 8194
use cut_M1M2_2x1 
transform 1 0 1060 0 1 16590
box 1060 16590 1244 16658
use cut_M1M2_2x1 
transform 1 0 4516 0 1 12354
box 4516 12354 4700 12422
use cut_M1M3_2x1 
transform 1 0 1060 0 1 20826
box 1060 20826 1260 20902
use cut_M1M3_2x1 
transform 1 0 4516 0 1 16590
box 4516 16590 4716 16666
use cut_M1M2_2x1 
transform 1 0 4516 0 1 20826
box 4516 20826 4700 20894
use cut_M2M4_2x1 
transform 1 0 5748 0 1 3124
box 5748 3124 5948 3200
use cut_M1M3_2x1 
transform 1 0 1060 0 1 3882
box 1060 3882 1260 3958
use cut_M3M4_2x1 
transform 1 0 5748 0 1 1204
box 5748 1204 5948 1280
use cut_M3M4_2x1 
transform 1 0 5748 0 1 2164
box 5748 2164 5948 2240
use cut_M1M4_1x2 
transform 1 0 39532 0 1 0
box 39532 0 39608 200
use cut_M1M4_1x2 
transform 1 0 39532 0 1 404
box 39532 404 39608 604
use cut_M1M4_1x2 
transform 1 0 39532 0 1 1364
box 39532 1364 39608 1564
use cut_M1M4_1x2 
transform 1 0 39532 0 1 2324
box 39532 2324 39608 2524
<< labels >>
flabel locali s 39532 0 39832 22068 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 4516 20826 5092 21046 0 FreeSans 400 0 0 0 VLPFZ
port 1 nsew
flabel locali s 1060 3882 1636 4102 0 FreeSans 400 0 0 0 VLPF
port 3 nsew
<< end >>
