magic
tech sky130B
magscale 1 2
timestamp 1679853665
<< locali >>
rect 0 5520 4056 5760
rect 0 240 240 5520
rect 384 5136 3672 5376
rect 384 624 624 5136
rect 1200 3026 1428 3086
rect 1368 2382 1428 3026
rect 1200 2322 1428 2382
rect 1368 1590 1428 2322
rect 1368 1530 1632 1590
rect 3432 624 3672 5136
rect 384 384 3672 624
rect 3816 240 4056 5520
rect 0 0 4056 240
<< metal1 >>
rect 1200 4786 1428 4846
rect 1368 4054 1428 4786
rect 1368 3994 1632 4054
rect 1092 3730 1200 3790
rect 972 3670 1152 3730
rect 972 3290 1032 3670
rect 1368 3438 1428 3994
rect 1200 3378 1428 3438
rect 1524 3290 1632 3350
rect 972 3230 1584 3290
rect 972 1326 1032 3230
rect 1200 2674 1428 2734
rect 1368 2470 1428 2674
rect 1368 2410 1632 2470
rect 972 1266 1200 1326
<< metal2 >>
rect 1632 4934 3948 4950
rect 1632 4874 4056 4934
rect 108 4142 1200 4158
rect 0 4082 1200 4142
rect 1632 2822 3948 2838
rect 1632 2762 4056 2822
rect 108 1678 1200 1694
rect 0 1618 1200 1678
<< metal3 >>
rect 1516 384 1732 4992
rect 2308 768 2524 5760
use cut_M1M2_2x1  cut_M1M2_2x1_0
timestamp 1677625200
transform 1 0 1124 0 1 3730
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_1
timestamp 1677625200
transform 1 0 1556 0 1 3290
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_2
timestamp 1677625200
transform 1 0 1124 0 1 1266
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_3
timestamp 1677625200
transform 1 0 1092 0 1 4786
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_4
timestamp 1677625200
transform 1 0 1524 0 1 3994
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_5
timestamp 1677625200
transform 1 0 1092 0 1 3378
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_6
timestamp 1677625200
transform 1 0 1524 0 1 2410
box 0 0 184 68
use cut_M1M2_2x1  cut_M1M2_2x1_7
timestamp 1677625200
transform 1 0 1092 0 1 2674
box 0 0 184 68
use cut_M1M3_2x1  cut_M1M3_2x1_0
timestamp 1677625200
transform 1 0 1524 0 1 4874
box 0 0 200 76
use cut_M1M3_2x1  cut_M1M3_2x1_1
timestamp 1677625200
transform 1 0 1524 0 1 2762
box 0 0 200 76
use cut_M1M3_2x1  cut_M1M3_2x1_2
timestamp 1677625200
transform 1 0 1108 0 1 4082
box 0 0 200 76
use cut_M1M3_2x1  cut_M1M3_2x1_3
timestamp 1677625200
transform 1 0 1108 0 1 1618
box 0 0 200 76
use cut_M1M4_2x1  cut_M1M4_2x1_0
timestamp 1677625200
transform 1 0 2316 0 1 5520
box 0 0 200 76
use cut_M1M4_2x1  cut_M1M4_2x1_1
timestamp 1677625200
transform 1 0 1524 0 1 384
box 0 0 200 76
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_TAPCELLB_CV#1  xa0 ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 0
transform 1 0 768 0 1 768
box 0 0 1 1
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFTSPCX1_CV  xa1 ../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1679853665
transform 1 0 768 0 1 1120
box -180 -132 2700 1188
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV#1  xa2 ../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1679853665
transform 1 0 768 0 1 2176
box -180 -132 2700 484
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV#1  xa2a
timestamp 1679853665
transform 1 0 768 0 1 2528
box -180 -132 2700 484
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_NRX1_CV  xa3 ../sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1679853665
transform 1 0 768 0 1 2880
box -180 -132 2700 836
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_DFTSPCX1_CV  xa5
timestamp 1679853665
transform 1 0 768 0 1 3584
box -180 -132 2700 1188
use ../../sun_tr_sky130nm/design/SUN_TR_SKY130NM/SUNTR_IVX1_CV#1  xa6
timestamp 1679853665
transform 1 0 768 0 1 4640
box -180 -132 2700 484
<< labels >>
flabel locali s 3432 384 3672 5376 0 FreeSans 400 0 0 0 AVSS
port 6 nsew
flabel locali s 3816 0 4056 5760 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel metal2 s 3840 2762 4056 2822 0 FreeSans 400 0 0 0 CP_UP_N
port 2 nsew
flabel metal2 s 0 1618 216 1678 0 FreeSans 400 0 0 0 CK_REF
port 3 nsew
flabel metal2 s 3840 4874 4056 4934 0 FreeSans 400 0 0 0 CP_DOWN
port 4 nsew
flabel metal2 s 0 4082 216 4142 0 FreeSans 400 0 0 0 CK_FB
port 5 nsew
<< end >>
