magic
tech sky130B
magscale 1 2
timestamp 1677625200
<< checkpaint >>
rect 0 0 56080 54840
<< locali >>
rect 55312 528 55552 54312
rect 528 528 55552 768
rect 528 54072 55552 54312
rect 528 528 768 54312
rect 55312 528 55552 54312
rect 55840 0 56080 54840
rect 0 0 56080 240
rect 0 54600 56080 54840
rect 0 0 240 54840
rect 55840 0 56080 54840
<< m2 >>
rect 1056 9138 1272 9198
rect 1056 2674 1272 2734
rect 1056 7730 1272 7790
<< m1 >>
rect 2580 39652 2796 39712
use SUN_PLL_PFD xaa0
transform 1 0 1056 0 1 1056
box 1056 1056 5112 6816
use SUN_PLL_CP xaa1
transform 1 0 1056 0 1 6816
box 1056 6816 5112 12752
use SUN_PLL_KICK xaa3
transform 1 0 1056 0 1 12752
box 1056 12752 5184 23264
use SUN_PLL_BUF xaa4
transform 1 0 1056 0 1 23264
box 1056 23264 15408 34304
use SUN_PLL_ROSC xaa5
transform 1 0 1056 0 1 34304
box 1056 34304 7632 39712
use SUN_PLL_DIVN xaa6
transform 1 0 1056 0 1 39712
box 1056 39712 15192 46748
use SUN_PLL_LPF xbb0
transform 1 0 15192 0 1 1056
box 15192 1056 55024 50904
use SUN_PLL_BIAS xbb1
transform 1 0 15192 0 1 50904
box 15192 50904 17220 53784
<< labels >>
flabel locali s 55312 528 55552 54312 0 FreeSans 400 0 0 0 AVSS
port 2 nsew
flabel locali s 55840 0 56080 54840 0 FreeSans 400 0 0 0 AVDD
port 1 nsew
flabel m2 s 1056 9138 1272 9198 0 FreeSans 400 0 0 0 PWRUP_1V8
port 3 nsew
flabel m2 s 1056 2674 1272 2734 0 FreeSans 400 0 0 0 CK_REF
port 4 nsew
flabel m1 s 2580 39652 2796 39712 0 FreeSans 400 0 0 0 CK
port 5 nsew
flabel m2 s 1056 7730 1272 7790 0 FreeSans 400 0 0 0 IBPSR_1U
port 6 nsew
<< end >>
