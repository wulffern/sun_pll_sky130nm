magic
tech sky130B
magscale 1 1
timestamp 1720908000
<< checkpaint >>
rect 0 0 38 100
<< locali >>
rect 0 0 34 92
<< m1 >>
rect 0 0 34 92
<< m2 >>
rect 0 0 38 100
<< m3 >>
rect 0 0 38 100
<< viali >>
rect 3 6 31 86
<< v1 >>
rect 3 6 31 86
<< v2 >>
rect 3 6 35 94
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 38 100
<< end >>
